/* Verilog model created from schematic Trying.sch -- Aug 14, 2020 14:52 */

module Trying;



load_register I2 ();

endmodule // Trying
