/* Verilog model created from schematic Top.sch -- Aug 13, 2020 20:32 */

module Top;




endmodule // Top
