// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.0.396.4
// Netlist written on Thu Aug 13 20:23:44 2020
//
// Verilog Description of module behave1p_mem
//

module behave1p_mem (d_out, wr_en, rd_en, clk, d_in, addr) /* synthesis syn_module_defined=1 */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(7[8:20])
    output [7:0]d_out;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(21[26:31])
    input wr_en;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(17[16:21])
    input rd_en;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(17[23:28])
    input clk;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(17[30:33])
    input [7:0]d_in;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(18[21:25])
    input [7:0]addr;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(19[27:31])
    
    wire clk_c /* synthesis is_clock=1, SET_AS_NETWORK=clk_c */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(17[30:33])
    
    wire n12909, wr_en_c, rd_en_c, d_in_c_7, d_in_c_6, d_in_c_5, 
        d_in_c_4, d_in_c_3, d_in_c_2, d_in_c_1, d_in_c_0, addr_c_7, 
        addr_c_6, addr_c_5, addr_c_4, addr_c_3, addr_c_2, addr_c_1, 
        addr_c_0, d_out_c_7, d_out_c_6, d_out_c_5, d_out_c_4, d_out_c_3, 
        d_out_c_2, d_out_c_1, d_out_c_0;
    wire [7:0]r_addr;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(23[21:27])
    wire [7:0]\array[0] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[1] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[2] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[3] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[4] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[5] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[6] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[7] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[8] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[9] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[10] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[11] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[12] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[13] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[14] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[15] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[16] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[17] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[18] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[19] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[20] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[21] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[22] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[23] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[24] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[25] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[26] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[27] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[28] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[29] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[30] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[31] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[32] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[33] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[34] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[35] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[36] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[37] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[38] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[39] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[40] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[41] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[42] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[43] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[44] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[45] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[46] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[47] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[48] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[49] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[50] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[51] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[52] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[53] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[54] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[55] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[56] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[57] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[58] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[59] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[60] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[61] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[62] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[63] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[64] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[65] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[66] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[67] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[68] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[69] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[70] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[71] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[72] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[73] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[74] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[75] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[76] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[77] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[78] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[79] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[80] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[81] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[82] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[83] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[84] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[85] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[86] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[87] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[88] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[89] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[90] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[91] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[92] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[93] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[94] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[95] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[96] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[97] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[98] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[99] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[100] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[101] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[102] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[103] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[104] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[105] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[106] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[107] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[108] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[109] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[110] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[111] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[112] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[113] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[114] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[115] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[116] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[117] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[118] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[119] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[120] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[121] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[122] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[123] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[124] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[125] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[126] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[127] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[128] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[129] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[130] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[131] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[132] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[133] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[134] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[135] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[136] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[137] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[138] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[139] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[140] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[141] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[142] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[143] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[144] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[145] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[146] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[147] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[148] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[149] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[150] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[151] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[152] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[153] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[154] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[155] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[156] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[157] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[158] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[159] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[160] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[161] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[162] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[163] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[164] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[165] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[166] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[167] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[168] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[169] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[170] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[171] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[172] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[173] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[174] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[175] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[176] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[177] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[178] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[179] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[180] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[181] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[182] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[183] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[184] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[185] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[186] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[187] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[188] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[189] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[190] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[191] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[192] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[193] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[194] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[195] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[196] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[197] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[198] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[199] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[200] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[201] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[202] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[203] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[204] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[205] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[206] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[207] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[208] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[209] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[210] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[211] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[212] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[213] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[214] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[215] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[216] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[217] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[218] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[219] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[220] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[221] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[222] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[223] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[224] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[225] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[226] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[227] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[228] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[229] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[230] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[231] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[232] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[233] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[234] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[235] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[236] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[237] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[238] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[239] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[240] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[241] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[242] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[243] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[244] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[245] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[246] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[247] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[248] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[249] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[250] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[251] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[252] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[253] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[254] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]\array[255] ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(25[30:35])
    wire [7:0]array_0__7__N_4097;
    wire [7:0]array_0__7__N_4089;
    wire [7:0]array_0__7__N_4081;
    wire [7:0]array_0__7__N_4073;
    wire [7:0]array_0__7__N_4065;
    wire [7:0]array_0__7__N_4057;
    wire [7:0]array_0__7__N_4049;
    wire [7:0]array_0__7__N_4041;
    wire [7:0]array_0__7__N_4033;
    wire [7:0]array_0__7__N_4025;
    wire [7:0]array_0__7__N_4017;
    wire [7:0]array_0__7__N_4009;
    wire [7:0]array_0__7__N_4001;
    wire [7:0]array_0__7__N_3993;
    wire [7:0]array_0__7__N_3985;
    wire [7:0]array_0__7__N_3977;
    wire [7:0]array_0__7__N_3969;
    wire [7:0]array_0__7__N_3961;
    wire [7:0]array_0__7__N_3953;
    wire [7:0]array_0__7__N_3945;
    wire [7:0]array_0__7__N_3937;
    wire [7:0]array_0__7__N_3929;
    wire [7:0]array_0__7__N_3921;
    wire [7:0]array_0__7__N_3913;
    wire [7:0]array_0__7__N_3905;
    wire [7:0]array_0__7__N_3897;
    wire [7:0]array_0__7__N_3889;
    wire [7:0]array_0__7__N_3881;
    wire [7:0]array_0__7__N_3873;
    wire [7:0]array_0__7__N_3865;
    wire [7:0]array_0__7__N_3857;
    wire [7:0]array_0__7__N_3849;
    wire [7:0]array_0__7__N_3841;
    wire [7:0]array_0__7__N_3833;
    wire [7:0]array_0__7__N_3825;
    wire [7:0]array_0__7__N_3817;
    wire [7:0]array_0__7__N_3809;
    wire [7:0]array_0__7__N_3801;
    wire [7:0]array_0__7__N_3793;
    wire [7:0]array_0__7__N_3785;
    wire [7:0]array_0__7__N_3777;
    wire [7:0]array_0__7__N_3769;
    wire [7:0]array_0__7__N_3761;
    wire [7:0]array_0__7__N_3753;
    wire [7:0]array_0__7__N_3745;
    wire [7:0]array_0__7__N_3737;
    wire [7:0]array_0__7__N_3729;
    wire [7:0]array_0__7__N_3721;
    wire [7:0]array_0__7__N_3713;
    wire [7:0]array_0__7__N_3705;
    wire [7:0]array_0__7__N_3697;
    wire [7:0]array_0__7__N_3689;
    wire [7:0]array_0__7__N_3681;
    wire [7:0]array_0__7__N_3673;
    wire [7:0]array_0__7__N_3665;
    wire [7:0]array_0__7__N_3657;
    wire [7:0]array_0__7__N_3649;
    wire [7:0]array_0__7__N_3641;
    wire [7:0]array_0__7__N_3633;
    wire [7:0]array_0__7__N_3625;
    wire [7:0]array_0__7__N_3617;
    wire [7:0]array_0__7__N_3609;
    wire [7:0]array_0__7__N_3601;
    wire [7:0]array_0__7__N_3593;
    wire [7:0]array_0__7__N_3585;
    wire [7:0]array_0__7__N_3577;
    wire [7:0]array_0__7__N_3569;
    wire [7:0]array_0__7__N_3561;
    wire [7:0]array_0__7__N_3553;
    wire [7:0]array_0__7__N_3545;
    wire [7:0]array_0__7__N_3537;
    wire [7:0]array_0__7__N_3529;
    wire [7:0]array_0__7__N_3521;
    wire [7:0]array_0__7__N_3513;
    wire [7:0]array_0__7__N_3505;
    wire [7:0]array_0__7__N_3497;
    wire [7:0]array_0__7__N_3489;
    wire [7:0]array_0__7__N_3481;
    wire [7:0]array_0__7__N_3473;
    wire [7:0]array_0__7__N_3465;
    wire [7:0]array_0__7__N_3457;
    wire [7:0]array_0__7__N_3449;
    wire [7:0]array_0__7__N_3441;
    wire [7:0]array_0__7__N_3433;
    wire [7:0]array_0__7__N_3425;
    wire [7:0]array_0__7__N_3417;
    wire [7:0]array_0__7__N_3409;
    wire [7:0]array_0__7__N_3401;
    wire [7:0]array_0__7__N_3393;
    wire [7:0]array_0__7__N_3385;
    wire [7:0]array_0__7__N_3377;
    wire [7:0]array_0__7__N_3369;
    wire [7:0]array_0__7__N_3361;
    wire [7:0]array_0__7__N_3353;
    wire [7:0]array_0__7__N_3345;
    wire [7:0]array_0__7__N_3337;
    wire [7:0]array_0__7__N_3329;
    wire [7:0]array_0__7__N_3321;
    wire [7:0]array_0__7__N_3313;
    wire [7:0]array_0__7__N_3305;
    wire [7:0]array_0__7__N_3297;
    wire [7:0]array_0__7__N_3289;
    wire [7:0]array_0__7__N_3281;
    wire [7:0]array_0__7__N_3273;
    wire [7:0]array_0__7__N_3265;
    wire [7:0]array_0__7__N_3257;
    wire [7:0]array_0__7__N_3249;
    wire [7:0]array_0__7__N_3241;
    wire [7:0]array_0__7__N_3233;
    wire [7:0]array_0__7__N_3225;
    wire [7:0]array_0__7__N_3217;
    wire [7:0]array_0__7__N_3209;
    wire [7:0]array_0__7__N_3201;
    wire [7:0]array_0__7__N_3193;
    wire [7:0]array_0__7__N_3185;
    wire [7:0]array_0__7__N_3177;
    wire [7:0]array_0__7__N_3169;
    wire [7:0]array_0__7__N_3161;
    wire [7:0]array_0__7__N_3153;
    wire [7:0]array_0__7__N_3145;
    wire [7:0]array_0__7__N_3137;
    wire [7:0]array_0__7__N_3129;
    wire [7:0]array_0__7__N_3121;
    wire [7:0]array_0__7__N_3113;
    wire [7:0]array_0__7__N_3105;
    wire [7:0]array_0__7__N_3097;
    wire [7:0]array_0__7__N_3089;
    wire [7:0]array_0__7__N_3081;
    wire [7:0]array_0__7__N_3073;
    wire [7:0]array_0__7__N_3065;
    wire [7:0]array_0__7__N_3057;
    wire [7:0]array_0__7__N_3049;
    wire [7:0]array_0__7__N_3041;
    wire [7:0]array_0__7__N_3033;
    wire [7:0]array_0__7__N_3025;
    wire [7:0]array_0__7__N_3017;
    wire [7:0]array_0__7__N_3009;
    wire [7:0]array_0__7__N_3001;
    wire [7:0]array_0__7__N_2993;
    wire [7:0]array_0__7__N_2985;
    wire [7:0]array_0__7__N_2977;
    wire [7:0]array_0__7__N_2969;
    wire [7:0]array_0__7__N_2961;
    wire [7:0]array_0__7__N_2953;
    wire [7:0]array_0__7__N_2945;
    wire [7:0]array_0__7__N_2937;
    wire [7:0]array_0__7__N_2929;
    wire [7:0]array_0__7__N_2921;
    wire [7:0]array_0__7__N_2913;
    wire [7:0]array_0__7__N_2905;
    wire [7:0]array_0__7__N_2897;
    wire [7:0]array_0__7__N_2889;
    wire [7:0]array_0__7__N_2881;
    wire [7:0]array_0__7__N_2873;
    wire [7:0]array_0__7__N_2865;
    wire [7:0]array_0__7__N_2857;
    wire [7:0]array_0__7__N_2849;
    wire [7:0]array_0__7__N_2841;
    wire [7:0]array_0__7__N_2833;
    wire [7:0]array_0__7__N_2825;
    wire [7:0]array_0__7__N_2817;
    wire [7:0]array_0__7__N_2809;
    wire [7:0]array_0__7__N_2801;
    wire [7:0]array_0__7__N_2793;
    wire [7:0]array_0__7__N_2785;
    wire [7:0]array_0__7__N_2777;
    wire [7:0]array_0__7__N_2769;
    wire [7:0]array_0__7__N_2761;
    wire [7:0]array_0__7__N_2753;
    wire [7:0]array_0__7__N_2745;
    wire [7:0]array_0__7__N_2737;
    wire [7:0]array_0__7__N_2729;
    wire [7:0]array_0__7__N_2721;
    wire [7:0]array_0__7__N_2713;
    wire [7:0]array_0__7__N_2705;
    wire [7:0]array_0__7__N_2697;
    wire [7:0]array_0__7__N_2689;
    wire [7:0]array_0__7__N_2681;
    wire [7:0]array_0__7__N_2673;
    wire [7:0]array_0__7__N_2665;
    wire [7:0]array_0__7__N_2657;
    wire [7:0]array_0__7__N_2649;
    wire [7:0]array_0__7__N_2641;
    wire [7:0]array_0__7__N_2633;
    wire [7:0]array_0__7__N_2625;
    wire [7:0]array_0__7__N_2617;
    wire [7:0]array_0__7__N_2609;
    wire [7:0]array_0__7__N_2601;
    wire [7:0]array_0__7__N_2593;
    wire [7:0]array_0__7__N_2585;
    wire [7:0]array_0__7__N_2577;
    wire [7:0]array_0__7__N_2569;
    wire [7:0]array_0__7__N_2561;
    wire [7:0]array_0__7__N_2553;
    wire [7:0]array_0__7__N_2545;
    wire [7:0]array_0__7__N_2537;
    wire [7:0]array_0__7__N_2529;
    wire [7:0]array_0__7__N_2521;
    wire [7:0]array_0__7__N_2513;
    wire [7:0]array_0__7__N_2505;
    wire [7:0]array_0__7__N_2497;
    wire [7:0]array_0__7__N_2489;
    wire [7:0]array_0__7__N_2481;
    wire [7:0]array_0__7__N_2473;
    wire [7:0]array_0__7__N_2465;
    wire [7:0]array_0__7__N_2457;
    wire [7:0]array_0__7__N_2449;
    wire [7:0]array_0__7__N_2441;
    wire [7:0]array_0__7__N_2433;
    wire [7:0]array_0__7__N_2425;
    wire [7:0]array_0__7__N_2417;
    wire [7:0]array_0__7__N_2409;
    wire [7:0]array_0__7__N_2401;
    wire [7:0]array_0__7__N_2393;
    wire [7:0]array_0__7__N_2385;
    wire [7:0]array_0__7__N_2377;
    wire [7:0]array_0__7__N_2369;
    wire [7:0]array_0__7__N_2361;
    wire [7:0]array_0__7__N_2353;
    wire [7:0]array_0__7__N_2345;
    wire [7:0]array_0__7__N_2337;
    wire [7:0]array_0__7__N_2329;
    wire [7:0]array_0__7__N_2321;
    wire [7:0]array_0__7__N_2313;
    wire [7:0]array_0__7__N_2305;
    wire [7:0]array_0__7__N_2297;
    wire [7:0]array_0__7__N_2289;
    wire [7:0]array_0__7__N_2281;
    wire [7:0]array_0__7__N_2273;
    wire [7:0]array_0__7__N_2265;
    wire [7:0]array_0__7__N_2257;
    wire [7:0]array_0__7__N_2249;
    wire [7:0]array_0__7__N_2241;
    wire [7:0]array_0__7__N_2233;
    wire [7:0]array_0__7__N_2225;
    wire [7:0]array_0__7__N_2217;
    wire [7:0]array_0__7__N_2209;
    wire [7:0]array_0__7__N_2201;
    wire [7:0]array_0__7__N_2193;
    wire [7:0]array_0__7__N_2185;
    wire [7:0]array_0__7__N_2177;
    wire [7:0]array_0__7__N_2169;
    wire [7:0]array_0__7__N_2161;
    wire [7:0]array_0__7__N_2153;
    wire [7:0]array_0__7__N_2145;
    wire [7:0]array_0__7__N_2137;
    wire [7:0]array_0__7__N_2129;
    wire [7:0]array_0__7__N_2121;
    wire [7:0]array_0__7__N_2113;
    wire [7:0]array_0__7__N_2105;
    wire [7:0]array_0__7__N_2097;
    wire [7:0]array_0__7__N_2089;
    wire [7:0]array_0__7__N_2081;
    wire [7:0]array_0__7__N_2073;
    wire [7:0]array_0__7__N_2065;
    wire [7:0]array_0__7__N_2057;
    
    wire VCC_net, clk_c_enable_2057, maxfan_replicated_net_23, clk_c_enable_2056, 
        clk_c_enable_2007, clk_c_enable_1007, n15023, n15022, n15021, 
        n15020, n15019, n15018, n15017, n15016, n15015, n15014, 
        n15013, n15012, n15011, n15010, n15009, n15008, n15007, 
        n15006, n15005, n15004, n15003, n15002, n15001, n15000, 
        n14999, n14998, n14997, n14996, n14995, n14994, n14993, 
        n14992, n13903, n13902, n14434, n13901, n13900, n14433, 
        n14700, n13899, n13898, n14431, n13897, n13896, n14430, 
        n14699, n14832, n13895, n13894, n14429, n13893, n13892, 
        n14428, n14698, n13890, n13889, n14427, n13888, n13887, 
        n14426, n14697, n14831, n14898, n13886, n13885, n14425, 
        n13884, n13883, n14424, n14696, n13882, n13881, n14423, 
        n13880, n13879, n14422, n14695, n14830, n13878, n13877, 
        n14421, n13876, n13875, n14420, n14694, n13874, n13873, 
        n14419, n13872, n13871, n14418, n14692, n14829, n14897, 
        n14931, n13870, n13869, n14417, n13868, n13867, n14416, 
        n14691, n13866, n13865, n14415, n13864, n13863, n14414, 
        n14690, n14828, n13862, n13861, n14413, n13859, n13858, 
        n14412, n14689, n13857, n13856, n14411, n13855, n13854, 
        n14410, n14688, n14827, n14896, n13853, n13852, n14409, 
        n13851, n13850, n14408, n14686, n13849, n13848, n14407, 
        n13847, n13846, n14406, n14685, n14826, n13845, n13844, 
        n14405, n13843, n13842, n14404, n14684, n13841, n13840, 
        n14403, n13839, n13838, n14402, n14683, n14825, n14895, 
        n14930, GND_net, n13837, n13836, n14400, n13835, n13834, 
        n14399, n14682, n13833, n13832, n14398, n13831, n13830, 
        n14397, n14681, n14824, n13828, n13827, n14396, n13826, 
        n13825, n14395, n14680, n13824, n13823, n14394, n13822, 
        n13821, n14393, n14679, n14823, n14894, n13820, n13819, 
        n14392, n13818, n13817, n14391, n14678, n13816, n13815, 
        n14390, n13814, n13813, n14389, n14677, n14822, n13812, 
        n13811, n14388, n13810, n13809, n14387, n14676, n13808, 
        n13807, n14386, n13806, n13805, n14385, n14675, n14821, 
        n14893, n14929, n13804, n13803, n14384, n13802, n13801, 
        n14383, n14674, n13800, n13799, n14382, n13797, n13796, 
        n14381, n14673, n14820, n13795, n13794, n14380, n13793, 
        n13792, n14379, n14672, n13791, n13790, n14378, n13789, 
        n13788, n14377, n14671, n14819, n14892, n13787, n13786, 
        n14376, n13785, n13784, n14375, n14670, n13783, n13782, 
        n14374, n13781, n13780, n14373, n14669, n14817, n13779, 
        n13778, n14372, n13777, n13776, n14371, n14668, n13775, 
        n13774, n14369, n13773, n13772, n14368, n14667, n14816, 
        n14891, n14928, n14947, n13771, n13770, n14367, n13769, 
        n13768, n14366, n14666, n13766, n13765, n14365, n13764, 
        n13763, n14364, n14665, n14815, n13762, n13761, n14363, 
        n13760, n13759, n14362, n14664, n13758, n13757, n14361, 
        n13756, n13755, n14360, n14663, n14814, n14890, n13754, 
        n13753, n14359, n13752, n13751, n14358, n14662, n13750, 
        n13749, n14357, n13748, n13747, n14356, n14661, n14813, 
        n13746, n13745, n14355, n13744, n13743, n14354, n14660, 
        n13742, n13741, n14353, n13740, n13739, n14352, n14659, 
        n14812, n14889, n14927, n13738, n13737, n14351, n13735, 
        n13734, n14350, n14658, n13733, n13732, n14349, n13731, 
        n13730, n14348, n14657, n14811, n13729, n13728, n14347, 
        n13727, n13726, n14346, n14655, n13725, n13724, n14345, 
        n13723, n13722, n14344, n14654, n14810, n14888, n13721, 
        n13720, n14343, n13719, n13718, n14342, n14653, n13717, 
        n13716, n14341, n13715, n13714, n14340, n14652, n14809, 
        n13713, n13712, n14338, n13711, n13710, n14337, n14651, 
        n13709, n13708, n14336, n13707, n13706, n14335, n14650, 
        n14808, n14887, n14926, n14946, n13704, n13703, n14334, 
        n13702, n13701, n14333, n14649, n13700, n13699, n14332, 
        n13698, n13697, n14331, n14648, n14807, n13696, n13695, 
        n14330, n13694, n13693, n14329, n14647, n13692, n13691, 
        n14328, n13690, n13689, n14327, n14646, n14806, n14886, 
        n13688, n13687, n14326, n13686, n13685, n14325, n14645, 
        n13684, n13683, n14324, n13682, n13681, n14323, n14644, 
        n14805, n13680, n13679, n14322, n13678, n13677, n14321, 
        n14643, n13676, n13675, n14320, n13674, n13672, n14319, 
        n14642, n14804, n14885, n14925, n13671, n13670, n14318, 
        n13669, n13668, n14317, n14641, n13666, n13665, n14316, 
        n13664, n13663, n14315, n14640, n14803, n13662, n13661, 
        n14314, n13660, n13659, n14313, n14639, n13658, n13657, 
        n14312, n13656, n13655, n14311, n14638, n14802, n14884, 
        n13654, n13653, n14310, n13652, n13651, n14309, n14637, 
        n13650, n13649, n14307, n13648, n13647, n14306, n14636, 
        n14801, n13646, n13645, n14305, n13644, n13643, n14304, 
        n14635, n13642, n13641, n14303, n13640, n13639, n14302, 
        n14634, n14800, n14883, n14924, n14945, n13638, n13637, 
        n14301, n13635, n13634, n14300, n14633, n13633, n13632, 
        n14299, n13631, n13630, n14298, n14632, n14799, n13629, 
        n13628, n14297, n13627, n13626, n14296, n14631, n13625, 
        n13624, n14295, n13623, n13622, n14294, n14630, n14798, 
        n14882, n13621, n13620, n14293, n13619, n13618, n14292, 
        n14629, n13617, n13616, n14291, n13615, n13614, n14290, 
        n14628, n14797, n13613, n13612, n14289, n13611, n13610, 
        n14288, n14627, n13609, n13608, n14287, n13607, n13606, 
        n14286, n14626, n14796, n14881, n14923, n13604, n13603, 
        n14285, n13602, n13601, n14284, n14624, n13600, n13599, 
        n14283, n13598, n13597, n14282, n14623, n14795, n13596, 
        n13595, n14281, n13594, n13593, n14280, n14622, n13592, 
        n13591, n14279, n13590, n13589, n14278, n14621, n14794, 
        n14879, n13588, n13587, n14276, n13586, n13585, n14275, 
        n14620, n13584, n13583, n14274, n13582, n13581, n14273, 
        n14619, n14793, n13580, n13579, n14272, n13578, n13577, 
        n14271, n14618, n13576, n13575, n14270, n13573, n13572, 
        n14269, n14617, n14792, n14878, n14922, n14944, n13571, 
        n13570, n14268, n13569, n13568, n14267, n14616, n13567, 
        n13566, n14266, n13565, n13564, n14265, n14615, n14791, 
        n13563, n13562, n14264, n13561, n13560, n14263, n14614, 
        n13559, n13558, n14262, n13557, n13556, n14261, n14613, 
        n14790, n14877, n13555, n13554, n14260, n13553, n13552, 
        n14259, n14612, n13551, n13550, n14258, n13549, n13548, 
        n14257, n14611, n14789, n13547, n13546, n14256, n13545, 
        n13544, n14255, n14610, n13542, n13541, n14254, n13540, 
        n13539, n14253, n14609, n14788, n14876, n14921, n13538, 
        n13537, n14252, n13536, n13535, n14251, n14608, n13534, 
        n13533, n14250, n13532, n13531, n14249, n14607, n14786, 
        n13530, n13529, n14248, n13528, n13527, n14247, n14606, 
        n13526, n13525, n14245, n13524, n13523, n14244, n14605, 
        n14785, n14875, n13522, n13521, n14243, n13520, n13519, 
        n14242, n14604, n13518, n13517, n14241, n13516, n13515, 
        n14240, n14603, n14784, n13514, n13513, n14239, n13511, 
        n13510, n14238, n14602, n13509, n13508, n14237, n13507, 
        n13506, n14236, n14601, n14783, n14874, n14920, n14943, 
        n13505, n13504, n14235, n13503, n13502, n14234, n14600, 
        n13501, n13500, n14233, n13499, n13498, n14232, n14599, 
        n14782, n13497, n13496, n14231, n13495, n13494, n14230, 
        n14598, n13493, n13492, n14229, n13491, n13490, n14228, 
        n14597, n14781, n14873, n13489, n13488, n14227, n13487, 
        n13486, n14226, n14596, n13485, n13484, n14225, n13483, 
        n13482, n14224, n14595, n14780, n13480, n13479, n14223, 
        n13478, n13477, n14222, n14593, n13476, n13475, n14221, 
        n13474, n13473, n14220, n14592, n14779, n14872, n14919, 
        n13472, n13471, n14219, n13470, n13469, n14218, n14591, 
        n13468, n13467, n14217, n13466, n13465, n14216, n14590, 
        n14778, n13464, n13463, n14214, n13462, n13461, n14213, 
        n14589, n13460, n13459, n14212, n13458, n13457, n14211, 
        n14588, n14777, n14871, n13456, n13455, n14210, n13454, 
        n13453, n14209, n14587, n13452, n13451, n14208, n13449, 
        n13448, n14207, n14586, n14776, n13447, n13446, n14206, 
        n13445, n13444, n14205, n14585, n13443, n13442, n14204, 
        n13441, n13440, n14203, n14584, n14775, n14870, n14918, 
        n14941, n13439, n13438, n14202, n13437, n13436, n14201, 
        n14583, n13435, n13434, n14200, n13433, n13432, n14199, 
        n14582, n14774, n13431, n13430, n14198, n13429, n13428, 
        n14197, n14581, n13427, n13426, n14196, n13425, n13424, 
        n14195, n14580, n14773, n14869, n13423, n13422, n14194, 
        n13421, n13420, n14193, n14579, n13419, n13417, n14192, 
        n13416, n13415, n14191, n14578, n14772, n13414, n13413, 
        n14190, n13411, n13410, n14189, n14577, n13409, n13408, 
        n14188, n13407, n13406, n14187, n14576, n14771, n14868, 
        n14917, n13405, n13404, n14186, n13403, n13402, n14185, 
        n14575, n13401, n13400, n14184, n13399, n13398, n14182, 
        n14574, n14770, n13397, n13396, n14181, n13395, n13394, 
        n14180, n14573, n13393, n13392, n14179, n13391, n13390, 
        n14178, n14572, n14769, n14867, n13389, n13388, n14176, 
        n13387, n13386, n14175, n14571, n13385, n13384, n14174, 
        n13383, n13382, n14173, n14570, n14768, n13380, n13379, 
        n14172, n13378, n13377, n14171, n14569, n13376, n13375, 
        n14170, n13374, n13373, n14169, n14568, n14767, n14866, 
        n14916, n14940, n13372, n13371, n14168, n13370, n13369, 
        n14167, n14567, n13368, n13367, n14166, n13366, n13365, 
        n14165, n14566, n14766, n13364, n13363, n14164, n13362, 
        n13361, n14163, n14565, n13360, n13359, n14162, n13358, 
        n13357, n14161, n14564, n14765, n14865, n13356, n13355, 
        n14160, n13354, n13353, n14159, n14562, n13352, n13351, 
        n14158, n13349, n13348, n14157, n14561, n14764, n13347, 
        n13346, n14156, n13345, n13344, n14155, n14560, n13343, 
        n13342, n14154, n13341, n13340, n14153, n14559, n14763, 
        n14864, n14915, n13339, n13338, n14152, n13337, n13336, 
        n14151, n14558, n13335, n13334, n14150, n13333, n13332, 
        n14149, n14557, n14762, n13331, n13330, n14148, n13329, 
        n13328, n14147, n14556, n13327, n13326, n14145, n13325, 
        n13324, n14144, n14555, n14761, n14863, n13323, n13322, 
        n14143, n13321, n13320, n14142, n14554, n13318, n13317, 
        n14141, n13316, n13315, n14140, n14553, n14760, n13314, 
        n13313, n14139, n13312, n13311, n14138, n14552, n13310, 
        n13309, n14137, n13308, n13307, n14136, n14551, n14759, 
        n14862, n14914, n14939, n13306, n13305, n14135, n13304, 
        n13303, n14134, n14550, n13302, n13301, n14133, n13300, 
        n13299, n14132, n14549, n14758, n13298, n13297, n14131, 
        n13296, n13295, n14130, n14548, n13294, n13293, n14129, 
        n13292, n13291, n14128, n14547, n14757, n14861, n13290, 
        n13289, n14127, n13287, n13286, n14126, n14546, n13285, 
        n13284, n14125, n13283, n13282, n14124, n14545, n14755, 
        n13281, n13280, n14123, n13279, n13278, n14122, n14544, 
        n13277, n13276, n14121, n13275, n13274, n14120, n14543, 
        n14754, n14860, n14913, n13273, n13272, n14119, n13271, 
        n13270, n14118, n14542, n13269, n13268, n14117, n13267, 
        n13266, n14116, n14541, n14753, n13265, n13264, n14114, 
        n13263, n13262, n14113, n14540, n13261, n13260, n14112, 
        n13259, n13258, n14111, n14539, n14752, n14859, n13256, 
        n13255, n14110, n13254, n13253, n14109, n14538, n13252, 
        n13251, n14108, n13250, n13249, n14107, n14537, n14751, 
        n13248, n13247, n14106, n13246, n13245, n14105, n14536, 
        n13244, n13243, n14104, n13242, n13241, n14103, n14535, 
        n14750, n14858, n14912, n14938, n13240, n13239, n14102, 
        n13238, n13237, n14101, n14534, n13236, n13235, n14100, 
        n13234, n13233, n14099, n14533, n14749, n13232, n13231, 
        n14098, n13230, n13229, n14097, n14531, n13228, n13227, 
        n14096, n13225, n13224, n14095, n14530, n14748, n14857, 
        n13223, n13222, n14094, n13221, n13220, n14093, n14529, 
        n13219, n13218, n14092, n13217, n13216, n14091, n14528, 
        n14747, n13215, n13214, n14090, n13213, n13212, n14089, 
        n14527, n13211, n13210, n14088, n13209, n13208, n14087, 
        n14526, n14746, n14856, n14910, n13207, n13206, n14086, 
        n13205, n13204, n14085, n14525, n13203, n13202, n14083, 
        n13201, n13200, n14082, n14524, n14745, n13199, n13198, 
        n14081, n13197, n13196, n14080, n14523, n13194, n13193, 
        n14079, n13192, n13191, n14078, n14522, n14744, n14855, 
        n13190, n13189, n14077, n13188, n13187, n14076, n14521, 
        n13186, n13185, n14075, n13184, n13183, n14074, n14520, 
        n14743, n13182, n13181, n14073, n13180, n13179, n14072, 
        n14519, n13178, n13177, n14071, n13176, n13175, n14070, 
        n14518, n14742, n14854, n14909, n14937, n13174, n13173, 
        n14069, n13172, n13171, n14068, n14517, n13170, n13169, 
        n14067, n13168, n13167, n14066, n14516, n14741, n13166, 
        n13165, n14065, n13164, n13162, n14064, n14515, n13161, 
        n13160, n14063, n13159, n13158, n14062, n14514, n14740, 
        n14853, n13156, n13155, n14061, n13154, n13153, n14060, 
        n14513, n13152, n13151, n14059, n13150, n13149, n14058, 
        n14512, n14739, n13148, n13147, n14057, n13146, n13145, 
        n14056, n14511, n13144, n13143, n14055, n13142, n13141, 
        n14054, n14510, n14738, n14852, n14908, n13140, n13132, 
        n14052, n13131, n13130, n14051, n14509, n14942, n13129, 
        n14050, n13128, n13127, n14049, n14508, n14737, n14911, 
        n13125, n14048, n13124, n13123, n14047, n14507, n14880, 
        n13122, n14046, n13121, n13120, n14045, n14506, n14736, 
        n14851, n14849, n13119, n14044, n13118, n13117, n14043, 
        n14505, n14818, n13116, n14042, n13115, n13114, n14041, 
        n14504, n14735, n14787, n13113, n14040, n13112, n13111, 
        n14039, n14503, n14756, n13110, n14038, n13109, n13108, 
        n14037, n14502, n14734, n14850, n14907, n14936, n14725, 
        n13107, n14036, n13106, n13105, n14035, n14500, n13139, 
        n13104, n14034, n13103, n13102, n14033, n14499, n14733, 
        n14687, n13101, n14032, n13100, n13099, n14031, n14498, 
        n14656, n13098, n14030, n13097, n13096, n14029, n14497, 
        n14732, n14848, n14625, n13094, n14028, n13093, n13092, 
        n14027, n14496, n14594, n13091, n14026, n13090, n13089, 
        n14025, n14495, n14731, n14563, n13088, n14024, n13087, 
        n13086, n14023, n14494, n14532, n13085, n14021, n13084, 
        n13083, n14020, n14493, n14730, n14847, n14906, n14501, 
        n13082, n14019, n13081, n13080, n14018, n14492, n14470, 
        n13079, n14017, n13078, n13077, n14016, n14491, n14729, 
        n13138, n13076, n14015, n13075, n13074, n14014, n14490, 
        n14432, n13073, n14013, n13072, n13071, n14012, n14489, 
        n14728, n14846, n14401, n13070, n14011, n13069, n13068, 
        n14010, n14488, n14370, n13067, n14009, n13066, n13065, 
        n14008, n14487, n14727, n14339, n13063, n14007, n13062, 
        n13061, n14006, n14486, n14308, n13060, n14005, n13059, 
        n13058, n14004, n14485, n14726, n14845, n14905, n14935, 
        n14277, n13057, n14003, n13056, n13055, n14002, n14484, 
        n14246, n13054, n14001, n13053, n13052, n14000, n14483, 
        n14724, n14215, n13051, n13999, n13050, n13049, n13998, 
        n14482, n13137, n13048, n13997, n13047, n13046, n13996, 
        n14481, n14723, n14844, n14177, n13045, n13995, n13044, 
        n13043, n13994, n14480, n14146, n13042, n13993, n13041, 
        n13040, n13992, n14479, n14722, n14115, n13039, n13990, 
        n13038, n13037, n13989, n14478, n14084, n13036, n13988, 
        n13035, n13034, n13987, n14477, n14721, n14843, n14904, 
        n14053, n13032, n13986, n13031, n13030, n13985, n14476, 
        n14022, n13029, n13984, n13028, n13027, n13983, n14475, 
        n14720, n13991, n13026, n13982, n13025, n13024, n13981, 
        n14474, n13960, n13023, n13980, n13022, n13021, n13979, 
        n14473, n14719, n14842, n13136, n13020, n13978, n13019, 
        n13018, n13977, n14472, n13922, n13017, n13976, n13016, 
        n13015, n13975, n14471, n14718, n13891, n13014, n13974, 
        n13013, n13012, n13973, n14469, n13860, n13011, n13972, 
        n13010, n13009, n13971, n14468, n14717, n14841, n14903, 
        n14934, n13829, n13008, n13970, n13007, n13006, n13969, 
        n14467, n13798, n13005, n13968, n13004, n13003, n13967, 
        n14466, n14716, n13767, n13001, n13966, n13000, n12999, 
        n13965, n14465, n13736, n12998, n13964, n12997, n12996, 
        n13963, n14464, n14715, n14840, n13705, n12995, n13962, 
        n12994, n12993, n13961, n14463, n13135, n12992, n13959, 
        n12991, n12990, n13958, n14462, n14714, n13667, n12989, 
        n13957, n12988, n12987, n13956, n14461, n13636, n12986, 
        n13955, n12985, n12984, n13954, n14460, n14713, n14839, 
        n14902, n13605, n12983, n13953, n12982, n12981, n13952, 
        n14459, n13574, n12980, n13951, n12979, n12978, n13950, 
        n14458, n14712, n13543, n12977, n13949, n12976, n12975, 
        n13948, n14457, n13512, n12974, n13947, n12973, n12972, 
        n13946, n14456, n14711, n14838, n13481, n12970, n13945, 
        n12969, n12968, n13944, n14455, n13450, n12967, n13943, 
        n12966, n12965, n13942, n14454, n14710, n13134, n12964, 
        n13941, n12963, n12962, n13940, n14453, n13412, n12961, 
        n13939, n12960, n12959, n13938, n14452, n14709, n14837, 
        n14901, n14933, n13381, n12958, n13937, n12957, n12956, 
        n13936, n14451, n13350, n12955, n13935, n12954, n12953, 
        n13934, n14450, n14708, n13319, n12952, n13933, n12951, 
        n12950, n13932, n14449, n13288, n12949, n13931, n12948, 
        n12947, n13930, n14448, n14707, n14836, n13257, n12946, 
        n13929, n12945, n12944, n13927, n14447, n13226, n12943, 
        n13926, n12942, n12941, n13925, n14446, n14706, n13195, 
        n12939, n13924, n12938, n12937, n13923, n14445, n13133, 
        n12936, n13921, n12935, n12934, n13920, n14444, n14705, 
        n14835, n14900, n13157, n12933, n13919, n12932, n12931, 
        n13918, n14443, n13126, n12930, n13917, n12929, n12928, 
        n13916, n14442, n14704, n13095, n12927, n13915, n12926, 
        n12925, n13914, n14441, n13064, n12924, n13913, n12923, 
        n12922, n13912, n14440, n14703, n14834, n13033, n12921, 
        n13911, n12920, n12919, n13910, n14439, n13002, n12918, 
        n13909, n12917, n12916, n13908, n14437, n14702, n12971, 
        n12915, n13907, n12914, n12913, n13906, n14436, n12940, 
        n12912, n13905, n12911, n12910, n13904, n14435, n14701, 
        n14833, n14899, n14932;
    
    LUT4 i5165_3_lut (.A(\array[36] [4]), .B(\array[37] [4]), .C(r_addr[0]), 
         .Z(n13707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5165_3_lut.init = 16'hcaca;
    LUT4 i5164_3_lut (.A(\array[34] [4]), .B(\array[35] [4]), .C(r_addr[0]), 
         .Z(n13706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5164_3_lut.init = 16'hcaca;
    LUT4 i5163_3_lut (.A(\array[32] [4]), .B(\array[33] [4]), .C(r_addr[0]), 
         .Z(n13705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5163_3_lut.init = 16'hcaca;
    LUT4 i6248_3_lut (.A(\array[102] [0]), .B(\array[103] [0]), .C(r_addr[0]), 
         .Z(n14790)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6248_3_lut.init = 16'hcaca;
    LUT4 i6247_3_lut (.A(\array[100] [0]), .B(\array[101] [0]), .C(r_addr[0]), 
         .Z(n14789)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6247_3_lut.init = 16'hcaca;
    LUT4 i6098_3_lut (.A(\array[222] [7]), .B(\array[223] [7]), .C(r_addr[0]), 
         .Z(n14640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6098_3_lut.init = 16'hcaca;
    LUT4 i6097_3_lut (.A(\array[220] [7]), .B(\array[221] [7]), .C(r_addr[0]), 
         .Z(n14639)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6097_3_lut.init = 16'hcaca;
    LUT4 i6246_3_lut (.A(\array[98] [0]), .B(\array[99] [0]), .C(r_addr[0]), 
         .Z(n14788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6246_3_lut.init = 16'hcaca;
    LUT4 i6245_3_lut (.A(\array[96] [0]), .B(\array[97] [0]), .C(r_addr[0]), 
         .Z(n14787)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6245_3_lut.init = 16'hcaca;
    LUT4 i6096_3_lut (.A(\array[218] [7]), .B(\array[219] [7]), .C(r_addr[0]), 
         .Z(n14638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6096_3_lut.init = 16'hcaca;
    LUT4 i6095_3_lut (.A(\array[216] [7]), .B(\array[217] [7]), .C(r_addr[0]), 
         .Z(n14637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6095_3_lut.init = 16'hcaca;
    LUT4 i6094_3_lut (.A(\array[214] [7]), .B(\array[215] [7]), .C(r_addr[0]), 
         .Z(n14636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6094_3_lut.init = 16'hcaca;
    LUT4 i6093_3_lut (.A(\array[212] [7]), .B(\array[213] [7]), .C(r_addr[0]), 
         .Z(n14635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6093_3_lut.init = 16'hcaca;
    LUT4 i6092_3_lut (.A(\array[210] [7]), .B(\array[211] [7]), .C(r_addr[0]), 
         .Z(n14634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6092_3_lut.init = 16'hcaca;
    LUT4 i6091_3_lut (.A(\array[208] [7]), .B(\array[209] [7]), .C(r_addr[0]), 
         .Z(n14633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6091_3_lut.init = 16'hcaca;
    LUT4 i5781_3_lut (.A(\array[158] [6]), .B(\array[159] [6]), .C(r_addr[0]), 
         .Z(n14323)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5781_3_lut.init = 16'hcaca;
    LUT4 i5780_3_lut (.A(\array[156] [6]), .B(\array[157] [6]), .C(r_addr[0]), 
         .Z(n14322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5780_3_lut.init = 16'hcaca;
    LUT4 i5147_3_lut (.A(\array[30] [4]), .B(\array[31] [4]), .C(r_addr[0]), 
         .Z(n13689)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5147_3_lut.init = 16'hcaca;
    LUT4 i5146_3_lut (.A(\array[28] [4]), .B(\array[29] [4]), .C(r_addr[0]), 
         .Z(n13688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5146_3_lut.init = 16'hcaca;
    LUT4 i5145_3_lut (.A(\array[26] [4]), .B(\array[27] [4]), .C(r_addr[0]), 
         .Z(n13687)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5145_3_lut.init = 16'hcaca;
    LUT4 i5144_3_lut (.A(\array[24] [4]), .B(\array[25] [4]), .C(r_addr[0]), 
         .Z(n13686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5144_3_lut.init = 16'hcaca;
    LUT4 i5779_3_lut (.A(\array[154] [6]), .B(\array[155] [6]), .C(r_addr[0]), 
         .Z(n14321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5779_3_lut.init = 16'hcaca;
    LUT4 i5778_3_lut (.A(\array[152] [6]), .B(\array[153] [6]), .C(r_addr[0]), 
         .Z(n14320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5778_3_lut.init = 16'hcaca;
    LUT4 i6090_3_lut (.A(\array[206] [7]), .B(\array[207] [7]), .C(r_addr[0]), 
         .Z(n14632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6090_3_lut.init = 16'hcaca;
    LUT4 i6089_3_lut (.A(\array[204] [7]), .B(\array[205] [7]), .C(r_addr[0]), 
         .Z(n14631)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6089_3_lut.init = 16'hcaca;
    LUT4 i5143_3_lut (.A(\array[22] [4]), .B(\array[23] [4]), .C(r_addr[0]), 
         .Z(n13685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5143_3_lut.init = 16'hcaca;
    LUT4 i5142_3_lut (.A(\array[20] [4]), .B(\array[21] [4]), .C(r_addr[0]), 
         .Z(n13684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5142_3_lut.init = 16'hcaca;
    LUT4 i5141_3_lut (.A(\array[18] [4]), .B(\array[19] [4]), .C(r_addr[0]), 
         .Z(n13683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5141_3_lut.init = 16'hcaca;
    LUT4 i5140_3_lut (.A(\array[16] [4]), .B(\array[17] [4]), .C(r_addr[0]), 
         .Z(n13682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5140_3_lut.init = 16'hcaca;
    LUT4 i5777_3_lut (.A(\array[150] [6]), .B(\array[151] [6]), .C(r_addr[0]), 
         .Z(n14319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5777_3_lut.init = 16'hcaca;
    LUT4 i5776_3_lut (.A(\array[148] [6]), .B(\array[149] [6]), .C(r_addr[0]), 
         .Z(n14318)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5776_3_lut.init = 16'hcaca;
    LUT4 i5139_3_lut (.A(\array[14] [4]), .B(\array[15] [4]), .C(r_addr[0]), 
         .Z(n13681)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5139_3_lut.init = 16'hcaca;
    LUT4 i5138_3_lut (.A(\array[12] [4]), .B(\array[13] [4]), .C(r_addr[0]), 
         .Z(n13680)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5138_3_lut.init = 16'hcaca;
    LUT4 i5137_3_lut (.A(\array[10] [4]), .B(\array[11] [4]), .C(r_addr[0]), 
         .Z(n13679)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5137_3_lut.init = 16'hcaca;
    LUT4 i5136_3_lut (.A(\array[8] [4]), .B(\array[9] [4]), .C(r_addr[0]), 
         .Z(n13678)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5136_3_lut.init = 16'hcaca;
    LUT4 i5775_3_lut (.A(\array[146] [6]), .B(\array[147] [6]), .C(r_addr[0]), 
         .Z(n14317)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5775_3_lut.init = 16'hcaca;
    LUT4 i5774_3_lut (.A(\array[144] [6]), .B(\array[145] [6]), .C(r_addr[0]), 
         .Z(n14316)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5774_3_lut.init = 16'hcaca;
    LUT4 i6088_3_lut (.A(\array[202] [7]), .B(\array[203] [7]), .C(r_addr[0]), 
         .Z(n14630)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6088_3_lut.init = 16'hcaca;
    LUT4 i6087_3_lut (.A(\array[200] [7]), .B(\array[201] [7]), .C(r_addr[0]), 
         .Z(n14629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6087_3_lut.init = 16'hcaca;
    LUT4 i5135_3_lut (.A(\array[6] [4]), .B(\array[7] [4]), .C(r_addr[0]), 
         .Z(n13677)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5135_3_lut.init = 16'hcaca;
    LUT4 i5134_3_lut (.A(\array[4] [4]), .B(\array[5] [4]), .C(r_addr[0]), 
         .Z(n13676)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5134_3_lut.init = 16'hcaca;
    LUT4 i5133_3_lut (.A(\array[2] [4]), .B(\array[3] [4]), .C(r_addr[0]), 
         .Z(n13675)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5133_3_lut.init = 16'hcaca;
    LUT4 i5132_3_lut (.A(\array[0] [4]), .B(\array[1] [4]), .C(r_addr[0]), 
         .Z(n13674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5132_3_lut.init = 16'hcaca;
    LUT4 i5773_3_lut (.A(\array[142] [6]), .B(\array[143] [6]), .C(r_addr[0]), 
         .Z(n14315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5773_3_lut.init = 16'hcaca;
    LUT4 i5772_3_lut (.A(\array[140] [6]), .B(\array[141] [6]), .C(r_addr[0]), 
         .Z(n14314)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5772_3_lut.init = 16'hcaca;
    LUT4 i5771_3_lut (.A(\array[138] [6]), .B(\array[139] [6]), .C(r_addr[0]), 
         .Z(n14313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5771_3_lut.init = 16'hcaca;
    LUT4 i5770_3_lut (.A(\array[136] [6]), .B(\array[137] [6]), .C(r_addr[0]), 
         .Z(n14312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5770_3_lut.init = 16'hcaca;
    LUT4 i6086_3_lut (.A(\array[198] [7]), .B(\array[199] [7]), .C(r_addr[0]), 
         .Z(n14628)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6086_3_lut.init = 16'hcaca;
    LUT4 i6085_3_lut (.A(\array[196] [7]), .B(\array[197] [7]), .C(r_addr[0]), 
         .Z(n14627)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6085_3_lut.init = 16'hcaca;
    LUT4 i5769_3_lut (.A(\array[134] [6]), .B(\array[135] [6]), .C(r_addr[0]), 
         .Z(n14311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5769_3_lut.init = 16'hcaca;
    LUT4 i5768_3_lut (.A(\array[132] [6]), .B(\array[133] [6]), .C(r_addr[0]), 
         .Z(n14310)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5768_3_lut.init = 16'hcaca;
    LUT4 i5767_3_lut (.A(\array[130] [6]), .B(\array[131] [6]), .C(r_addr[0]), 
         .Z(n14309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5767_3_lut.init = 16'hcaca;
    LUT4 i5766_3_lut (.A(\array[128] [6]), .B(\array[129] [6]), .C(r_addr[0]), 
         .Z(n14308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5766_3_lut.init = 16'hcaca;
    LUT4 i6084_3_lut (.A(\array[194] [7]), .B(\array[195] [7]), .C(r_addr[0]), 
         .Z(n14626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6084_3_lut.init = 16'hcaca;
    LUT4 i6083_3_lut (.A(\array[192] [7]), .B(\array[193] [7]), .C(r_addr[0]), 
         .Z(n14625)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6083_3_lut.init = 16'hcaca;
    LUT4 i5109_3_lut (.A(\array[254] [3]), .B(\array[255] [3]), .C(r_addr[0]), 
         .Z(n13651)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5109_3_lut.init = 16'hcaca;
    LUT4 i5108_3_lut (.A(\array[252] [3]), .B(\array[253] [3]), .C(r_addr[0]), 
         .Z(n13650)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5108_3_lut.init = 16'hcaca;
    LUT4 i5107_3_lut (.A(\array[250] [3]), .B(\array[251] [3]), .C(r_addr[0]), 
         .Z(n13649)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5107_3_lut.init = 16'hcaca;
    LUT4 i5106_3_lut (.A(\array[248] [3]), .B(\array[249] [3]), .C(r_addr[0]), 
         .Z(n13648)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5106_3_lut.init = 16'hcaca;
    LUT4 i5105_3_lut (.A(\array[246] [3]), .B(\array[247] [3]), .C(r_addr[0]), 
         .Z(n13647)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5105_3_lut.init = 16'hcaca;
    LUT4 i5104_3_lut (.A(\array[244] [3]), .B(\array[245] [3]), .C(r_addr[0]), 
         .Z(n13646)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5104_3_lut.init = 16'hcaca;
    LUT4 i5103_3_lut (.A(\array[242] [3]), .B(\array[243] [3]), .C(r_addr[0]), 
         .Z(n13645)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5103_3_lut.init = 16'hcaca;
    LUT4 i5102_3_lut (.A(\array[240] [3]), .B(\array[241] [3]), .C(r_addr[0]), 
         .Z(n13644)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5102_3_lut.init = 16'hcaca;
    LUT4 i5101_3_lut (.A(\array[238] [3]), .B(\array[239] [3]), .C(r_addr[0]), 
         .Z(n13643)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5101_3_lut.init = 16'hcaca;
    LUT4 i5100_3_lut (.A(\array[236] [3]), .B(\array[237] [3]), .C(r_addr[0]), 
         .Z(n13642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5100_3_lut.init = 16'hcaca;
    LUT4 i5099_3_lut (.A(\array[234] [3]), .B(\array[235] [3]), .C(r_addr[0]), 
         .Z(n13641)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5099_3_lut.init = 16'hcaca;
    LUT4 i5098_3_lut (.A(\array[232] [3]), .B(\array[233] [3]), .C(r_addr[0]), 
         .Z(n13640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5098_3_lut.init = 16'hcaca;
    LUT4 i5097_3_lut (.A(\array[230] [3]), .B(\array[231] [3]), .C(r_addr[0]), 
         .Z(n13639)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5097_3_lut.init = 16'hcaca;
    LUT4 i5096_3_lut (.A(\array[228] [3]), .B(\array[229] [3]), .C(r_addr[0]), 
         .Z(n13638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5096_3_lut.init = 16'hcaca;
    LUT4 i5095_3_lut (.A(\array[226] [3]), .B(\array[227] [3]), .C(r_addr[0]), 
         .Z(n13637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5095_3_lut.init = 16'hcaca;
    LUT4 i5094_3_lut (.A(\array[224] [3]), .B(\array[225] [3]), .C(r_addr[0]), 
         .Z(n13636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5094_3_lut.init = 16'hcaca;
    LUT4 i5750_3_lut (.A(\array[126] [6]), .B(\array[127] [6]), .C(r_addr[0]), 
         .Z(n14292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5750_3_lut.init = 16'hcaca;
    LUT4 i5749_3_lut (.A(\array[124] [6]), .B(\array[125] [6]), .C(r_addr[0]), 
         .Z(n14291)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5749_3_lut.init = 16'hcaca;
    LUT4 i5748_3_lut (.A(\array[122] [6]), .B(\array[123] [6]), .C(r_addr[0]), 
         .Z(n14290)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5748_3_lut.init = 16'hcaca;
    LUT4 i5747_3_lut (.A(\array[120] [6]), .B(\array[121] [6]), .C(r_addr[0]), 
         .Z(n14289)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5747_3_lut.init = 16'hcaca;
    LUT4 i5746_3_lut (.A(\array[118] [6]), .B(\array[119] [6]), .C(r_addr[0]), 
         .Z(n14288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5746_3_lut.init = 16'hcaca;
    LUT4 i5745_3_lut (.A(\array[116] [6]), .B(\array[117] [6]), .C(r_addr[0]), 
         .Z(n14287)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5745_3_lut.init = 16'hcaca;
    LUT4 i5744_3_lut (.A(\array[114] [6]), .B(\array[115] [6]), .C(r_addr[0]), 
         .Z(n14286)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5744_3_lut.init = 16'hcaca;
    LUT4 i5743_3_lut (.A(\array[112] [6]), .B(\array[113] [6]), .C(r_addr[0]), 
         .Z(n14285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5743_3_lut.init = 16'hcaca;
    LUT4 i5742_3_lut (.A(\array[110] [6]), .B(\array[111] [6]), .C(r_addr[0]), 
         .Z(n14284)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5742_3_lut.init = 16'hcaca;
    LUT4 i5741_3_lut (.A(\array[108] [6]), .B(\array[109] [6]), .C(r_addr[0]), 
         .Z(n14283)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5741_3_lut.init = 16'hcaca;
    LUT4 i5078_3_lut (.A(\array[222] [3]), .B(\array[223] [3]), .C(r_addr[0]), 
         .Z(n13620)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5078_3_lut.init = 16'hcaca;
    LUT4 i5077_3_lut (.A(\array[220] [3]), .B(\array[221] [3]), .C(r_addr[0]), 
         .Z(n13619)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5077_3_lut.init = 16'hcaca;
    LUT4 i5076_3_lut (.A(\array[218] [3]), .B(\array[219] [3]), .C(r_addr[0]), 
         .Z(n13618)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5076_3_lut.init = 16'hcaca;
    LUT4 i5075_3_lut (.A(\array[216] [3]), .B(\array[217] [3]), .C(r_addr[0]), 
         .Z(n13617)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5075_3_lut.init = 16'hcaca;
    LUT4 i5740_3_lut (.A(\array[106] [6]), .B(\array[107] [6]), .C(r_addr[0]), 
         .Z(n14282)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5740_3_lut.init = 16'hcaca;
    LUT4 i5739_3_lut (.A(\array[104] [6]), .B(\array[105] [6]), .C(r_addr[0]), 
         .Z(n14281)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5739_3_lut.init = 16'hcaca;
    LUT4 i5074_3_lut (.A(\array[214] [3]), .B(\array[215] [3]), .C(r_addr[0]), 
         .Z(n13616)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5074_3_lut.init = 16'hcaca;
    LUT4 i5073_3_lut (.A(\array[212] [3]), .B(\array[213] [3]), .C(r_addr[0]), 
         .Z(n13615)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5073_3_lut.init = 16'hcaca;
    LUT4 i5072_3_lut (.A(\array[210] [3]), .B(\array[211] [3]), .C(r_addr[0]), 
         .Z(n13614)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5072_3_lut.init = 16'hcaca;
    LUT4 i5071_3_lut (.A(\array[208] [3]), .B(\array[209] [3]), .C(r_addr[0]), 
         .Z(n13613)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5071_3_lut.init = 16'hcaca;
    LUT4 i5738_3_lut (.A(\array[102] [6]), .B(\array[103] [6]), .C(r_addr[0]), 
         .Z(n14280)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5738_3_lut.init = 16'hcaca;
    LUT4 i5737_3_lut (.A(\array[100] [6]), .B(\array[101] [6]), .C(r_addr[0]), 
         .Z(n14279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5737_3_lut.init = 16'hcaca;
    LUT4 i5070_3_lut (.A(\array[206] [3]), .B(\array[207] [3]), .C(r_addr[0]), 
         .Z(n13612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5070_3_lut.init = 16'hcaca;
    LUT4 i5069_3_lut (.A(\array[204] [3]), .B(\array[205] [3]), .C(r_addr[0]), 
         .Z(n13611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5069_3_lut.init = 16'hcaca;
    LUT4 i5068_3_lut (.A(\array[202] [3]), .B(\array[203] [3]), .C(r_addr[0]), 
         .Z(n13610)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5068_3_lut.init = 16'hcaca;
    LUT4 i5067_3_lut (.A(\array[200] [3]), .B(\array[201] [3]), .C(r_addr[0]), 
         .Z(n13609)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5067_3_lut.init = 16'hcaca;
    LUT4 i5736_3_lut (.A(\array[98] [6]), .B(\array[99] [6]), .C(r_addr[0]), 
         .Z(n14278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5736_3_lut.init = 16'hcaca;
    LUT4 i5735_3_lut (.A(\array[96] [6]), .B(\array[97] [6]), .C(r_addr[0]), 
         .Z(n14277)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5735_3_lut.init = 16'hcaca;
    LUT4 i5066_3_lut (.A(\array[198] [3]), .B(\array[199] [3]), .C(r_addr[0]), 
         .Z(n13608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5066_3_lut.init = 16'hcaca;
    LUT4 i5065_3_lut (.A(\array[196] [3]), .B(\array[197] [3]), .C(r_addr[0]), 
         .Z(n13607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5065_3_lut.init = 16'hcaca;
    LUT4 i5064_3_lut (.A(\array[194] [3]), .B(\array[195] [3]), .C(r_addr[0]), 
         .Z(n13606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5064_3_lut.init = 16'hcaca;
    LUT4 i5063_3_lut (.A(\array[192] [3]), .B(\array[193] [3]), .C(r_addr[0]), 
         .Z(n13605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5063_3_lut.init = 16'hcaca;
    LUT4 i5047_3_lut (.A(\array[190] [3]), .B(\array[191] [3]), .C(r_addr[0]), 
         .Z(n13589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5047_3_lut.init = 16'hcaca;
    LUT4 i5046_3_lut (.A(\array[188] [3]), .B(\array[189] [3]), .C(r_addr[0]), 
         .Z(n13588)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5046_3_lut.init = 16'hcaca;
    LUT4 i5045_3_lut (.A(\array[186] [3]), .B(\array[187] [3]), .C(r_addr[0]), 
         .Z(n13587)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5045_3_lut.init = 16'hcaca;
    LUT4 i5044_3_lut (.A(\array[184] [3]), .B(\array[185] [3]), .C(r_addr[0]), 
         .Z(n13586)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5044_3_lut.init = 16'hcaca;
    LUT4 i5043_3_lut (.A(\array[182] [3]), .B(\array[183] [3]), .C(r_addr[0]), 
         .Z(n13585)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5043_3_lut.init = 16'hcaca;
    LUT4 i5042_3_lut (.A(\array[180] [3]), .B(\array[181] [3]), .C(r_addr[0]), 
         .Z(n13584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5042_3_lut.init = 16'hcaca;
    LUT4 i5041_3_lut (.A(\array[178] [3]), .B(\array[179] [3]), .C(r_addr[0]), 
         .Z(n13583)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5041_3_lut.init = 16'hcaca;
    LUT4 i5040_3_lut (.A(\array[176] [3]), .B(\array[177] [3]), .C(r_addr[0]), 
         .Z(n13582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5040_3_lut.init = 16'hcaca;
    LUT4 i5039_3_lut (.A(\array[174] [3]), .B(\array[175] [3]), .C(r_addr[0]), 
         .Z(n13581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5039_3_lut.init = 16'hcaca;
    LUT4 i5038_3_lut (.A(\array[172] [3]), .B(\array[173] [3]), .C(r_addr[0]), 
         .Z(n13580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5038_3_lut.init = 16'hcaca;
    LUT4 i5037_3_lut (.A(\array[170] [3]), .B(\array[171] [3]), .C(r_addr[0]), 
         .Z(n13579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5037_3_lut.init = 16'hcaca;
    LUT4 i5036_3_lut (.A(\array[168] [3]), .B(\array[169] [3]), .C(r_addr[0]), 
         .Z(n13578)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5036_3_lut.init = 16'hcaca;
    LUT4 i5035_3_lut (.A(\array[166] [3]), .B(\array[167] [3]), .C(r_addr[0]), 
         .Z(n13577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5035_3_lut.init = 16'hcaca;
    LUT4 i5034_3_lut (.A(\array[164] [3]), .B(\array[165] [3]), .C(r_addr[0]), 
         .Z(n13576)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5034_3_lut.init = 16'hcaca;
    LUT4 i5033_3_lut (.A(\array[162] [3]), .B(\array[163] [3]), .C(r_addr[0]), 
         .Z(n13575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5033_3_lut.init = 16'hcaca;
    LUT4 i5032_3_lut (.A(\array[160] [3]), .B(\array[161] [3]), .C(r_addr[0]), 
         .Z(n13574)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5032_3_lut.init = 16'hcaca;
    LUT4 i6067_3_lut (.A(\array[190] [7]), .B(\array[191] [7]), .C(r_addr[0]), 
         .Z(n14609)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6067_3_lut.init = 16'hcaca;
    LUT4 i6066_3_lut (.A(\array[188] [7]), .B(\array[189] [7]), .C(r_addr[0]), 
         .Z(n14608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6066_3_lut.init = 16'hcaca;
    LUT4 i6065_3_lut (.A(\array[186] [7]), .B(\array[187] [7]), .C(r_addr[0]), 
         .Z(n14607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6065_3_lut.init = 16'hcaca;
    LUT4 i6064_3_lut (.A(\array[184] [7]), .B(\array[185] [7]), .C(r_addr[0]), 
         .Z(n14606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6064_3_lut.init = 16'hcaca;
    LUT4 i6063_3_lut (.A(\array[182] [7]), .B(\array[183] [7]), .C(r_addr[0]), 
         .Z(n14605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6063_3_lut.init = 16'hcaca;
    LUT4 i6062_3_lut (.A(\array[180] [7]), .B(\array[181] [7]), .C(r_addr[0]), 
         .Z(n14604)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6062_3_lut.init = 16'hcaca;
    LUT4 i6322_3_lut (.A(\array[190] [0]), .B(\array[191] [0]), .C(r_addr[0]), 
         .Z(n14864)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6322_3_lut.init = 16'hcaca;
    LUT4 i6321_3_lut (.A(\array[188] [0]), .B(\array[189] [0]), .C(r_addr[0]), 
         .Z(n14863)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6321_3_lut.init = 16'hcaca;
    LUT4 i6061_3_lut (.A(\array[178] [7]), .B(\array[179] [7]), .C(r_addr[0]), 
         .Z(n14603)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6061_3_lut.init = 16'hcaca;
    LUT4 i6060_3_lut (.A(\array[176] [7]), .B(\array[177] [7]), .C(r_addr[0]), 
         .Z(n14602)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6060_3_lut.init = 16'hcaca;
    LUT4 i5719_3_lut (.A(\array[94] [6]), .B(\array[95] [6]), .C(r_addr[0]), 
         .Z(n14261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5719_3_lut.init = 16'hcaca;
    LUT4 i5718_3_lut (.A(\array[92] [6]), .B(\array[93] [6]), .C(r_addr[0]), 
         .Z(n14260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5718_3_lut.init = 16'hcaca;
    LUT4 i5717_3_lut (.A(\array[90] [6]), .B(\array[91] [6]), .C(r_addr[0]), 
         .Z(n14259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5717_3_lut.init = 16'hcaca;
    LUT4 i5716_3_lut (.A(\array[88] [6]), .B(\array[89] [6]), .C(r_addr[0]), 
         .Z(n14258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5716_3_lut.init = 16'hcaca;
    LUT4 i6059_3_lut (.A(\array[174] [7]), .B(\array[175] [7]), .C(r_addr[0]), 
         .Z(n14601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6059_3_lut.init = 16'hcaca;
    LUT4 i6058_3_lut (.A(\array[172] [7]), .B(\array[173] [7]), .C(r_addr[0]), 
         .Z(n14600)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6058_3_lut.init = 16'hcaca;
    LUT4 i5715_3_lut (.A(\array[86] [6]), .B(\array[87] [6]), .C(r_addr[0]), 
         .Z(n14257)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5715_3_lut.init = 16'hcaca;
    LUT4 i5714_3_lut (.A(\array[84] [6]), .B(\array[85] [6]), .C(r_addr[0]), 
         .Z(n14256)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5714_3_lut.init = 16'hcaca;
    LUT4 i5713_3_lut (.A(\array[82] [6]), .B(\array[83] [6]), .C(r_addr[0]), 
         .Z(n14255)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5713_3_lut.init = 16'hcaca;
    LUT4 i5712_3_lut (.A(\array[80] [6]), .B(\array[81] [6]), .C(r_addr[0]), 
         .Z(n14254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5712_3_lut.init = 16'hcaca;
    LUT4 i6057_3_lut (.A(\array[170] [7]), .B(\array[171] [7]), .C(r_addr[0]), 
         .Z(n14599)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6057_3_lut.init = 16'hcaca;
    LUT4 i6056_3_lut (.A(\array[168] [7]), .B(\array[169] [7]), .C(r_addr[0]), 
         .Z(n14598)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6056_3_lut.init = 16'hcaca;
    LUT4 i5711_3_lut (.A(\array[78] [6]), .B(\array[79] [6]), .C(r_addr[0]), 
         .Z(n14253)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5711_3_lut.init = 16'hcaca;
    LUT4 i5710_3_lut (.A(\array[76] [6]), .B(\array[77] [6]), .C(r_addr[0]), 
         .Z(n14252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5710_3_lut.init = 16'hcaca;
    LUT4 i5016_3_lut (.A(\array[158] [3]), .B(\array[159] [3]), .C(r_addr[0]), 
         .Z(n13558)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5016_3_lut.init = 16'hcaca;
    LUT4 i5015_3_lut (.A(\array[156] [3]), .B(\array[157] [3]), .C(r_addr[0]), 
         .Z(n13557)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5015_3_lut.init = 16'hcaca;
    LUT4 i5014_3_lut (.A(\array[154] [3]), .B(\array[155] [3]), .C(r_addr[0]), 
         .Z(n13556)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5014_3_lut.init = 16'hcaca;
    LUT4 i5013_3_lut (.A(\array[152] [3]), .B(\array[153] [3]), .C(r_addr[0]), 
         .Z(n13555)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5013_3_lut.init = 16'hcaca;
    LUT4 i5709_3_lut (.A(\array[74] [6]), .B(\array[75] [6]), .C(r_addr[0]), 
         .Z(n14251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5709_3_lut.init = 16'hcaca;
    LUT4 i5708_3_lut (.A(\array[72] [6]), .B(\array[73] [6]), .C(r_addr[0]), 
         .Z(n14250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5708_3_lut.init = 16'hcaca;
    LUT4 i6055_3_lut (.A(\array[166] [7]), .B(\array[167] [7]), .C(r_addr[0]), 
         .Z(n14597)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6055_3_lut.init = 16'hcaca;
    LUT4 i6054_3_lut (.A(\array[164] [7]), .B(\array[165] [7]), .C(r_addr[0]), 
         .Z(n14596)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6054_3_lut.init = 16'hcaca;
    LUT4 i6320_3_lut (.A(\array[186] [0]), .B(\array[187] [0]), .C(r_addr[0]), 
         .Z(n14862)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6320_3_lut.init = 16'hcaca;
    LUT4 i6319_3_lut (.A(\array[184] [0]), .B(\array[185] [0]), .C(r_addr[0]), 
         .Z(n14861)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6319_3_lut.init = 16'hcaca;
    LUT4 i5012_3_lut (.A(\array[150] [3]), .B(\array[151] [3]), .C(r_addr[0]), 
         .Z(n13554)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5012_3_lut.init = 16'hcaca;
    LUT4 i5011_3_lut (.A(\array[148] [3]), .B(\array[149] [3]), .C(r_addr[0]), 
         .Z(n13553)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5011_3_lut.init = 16'hcaca;
    LUT4 i5010_3_lut (.A(\array[146] [3]), .B(\array[147] [3]), .C(r_addr[0]), 
         .Z(n13552)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5010_3_lut.init = 16'hcaca;
    LUT4 i5009_3_lut (.A(\array[144] [3]), .B(\array[145] [3]), .C(r_addr[0]), 
         .Z(n13551)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5009_3_lut.init = 16'hcaca;
    LUT4 i5707_3_lut (.A(\array[70] [6]), .B(\array[71] [6]), .C(r_addr[0]), 
         .Z(n14249)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5707_3_lut.init = 16'hcaca;
    LUT4 i5706_3_lut (.A(\array[68] [6]), .B(\array[69] [6]), .C(r_addr[0]), 
         .Z(n14248)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5706_3_lut.init = 16'hcaca;
    LUT4 i5008_3_lut (.A(\array[142] [3]), .B(\array[143] [3]), .C(r_addr[0]), 
         .Z(n13550)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5008_3_lut.init = 16'hcaca;
    LUT4 i5007_3_lut (.A(\array[140] [3]), .B(\array[141] [3]), .C(r_addr[0]), 
         .Z(n13549)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5007_3_lut.init = 16'hcaca;
    LUT4 i5006_3_lut (.A(\array[138] [3]), .B(\array[139] [3]), .C(r_addr[0]), 
         .Z(n13548)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5006_3_lut.init = 16'hcaca;
    LUT4 i5005_3_lut (.A(\array[136] [3]), .B(\array[137] [3]), .C(r_addr[0]), 
         .Z(n13547)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5005_3_lut.init = 16'hcaca;
    LUT4 i5705_3_lut (.A(\array[66] [6]), .B(\array[67] [6]), .C(r_addr[0]), 
         .Z(n14247)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5705_3_lut.init = 16'hcaca;
    LUT4 i5704_3_lut (.A(\array[64] [6]), .B(\array[65] [6]), .C(r_addr[0]), 
         .Z(n14246)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5704_3_lut.init = 16'hcaca;
    LUT4 i6053_3_lut (.A(\array[162] [7]), .B(\array[163] [7]), .C(r_addr[0]), 
         .Z(n14595)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6053_3_lut.init = 16'hcaca;
    LUT4 i6052_3_lut (.A(\array[160] [7]), .B(\array[161] [7]), .C(r_addr[0]), 
         .Z(n14594)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6052_3_lut.init = 16'hcaca;
    LUT4 i5004_3_lut (.A(\array[134] [3]), .B(\array[135] [3]), .C(r_addr[0]), 
         .Z(n13546)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5004_3_lut.init = 16'hcaca;
    LUT4 i5003_3_lut (.A(\array[132] [3]), .B(\array[133] [3]), .C(r_addr[0]), 
         .Z(n13545)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5003_3_lut.init = 16'hcaca;
    LUT4 i5002_3_lut (.A(\array[130] [3]), .B(\array[131] [3]), .C(r_addr[0]), 
         .Z(n13544)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5002_3_lut.init = 16'hcaca;
    LUT4 i5001_3_lut (.A(\array[128] [3]), .B(\array[129] [3]), .C(r_addr[0]), 
         .Z(n13543)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5001_3_lut.init = 16'hcaca;
    LUT4 i6318_3_lut (.A(\array[182] [0]), .B(\array[183] [0]), .C(r_addr[0]), 
         .Z(n14860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6318_3_lut.init = 16'hcaca;
    LUT4 i6317_3_lut (.A(\array[180] [0]), .B(\array[181] [0]), .C(r_addr[0]), 
         .Z(n14859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6317_3_lut.init = 16'hcaca;
    LUT4 i4985_3_lut (.A(\array[126] [3]), .B(\array[127] [3]), .C(r_addr[0]), 
         .Z(n13527)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4985_3_lut.init = 16'hcaca;
    LUT4 i4984_3_lut (.A(\array[124] [3]), .B(\array[125] [3]), .C(r_addr[0]), 
         .Z(n13526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4984_3_lut.init = 16'hcaca;
    LUT4 i4983_3_lut (.A(\array[122] [3]), .B(\array[123] [3]), .C(r_addr[0]), 
         .Z(n13525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4983_3_lut.init = 16'hcaca;
    LUT4 i4982_3_lut (.A(\array[120] [3]), .B(\array[121] [3]), .C(r_addr[0]), 
         .Z(n13524)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4982_3_lut.init = 16'hcaca;
    LUT4 i4981_3_lut (.A(\array[118] [3]), .B(\array[119] [3]), .C(r_addr[0]), 
         .Z(n13523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4981_3_lut.init = 16'hcaca;
    LUT4 i4980_3_lut (.A(\array[116] [3]), .B(\array[117] [3]), .C(r_addr[0]), 
         .Z(n13522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4980_3_lut.init = 16'hcaca;
    LUT4 i4979_3_lut (.A(\array[114] [3]), .B(\array[115] [3]), .C(r_addr[0]), 
         .Z(n13521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4979_3_lut.init = 16'hcaca;
    LUT4 i4978_3_lut (.A(\array[112] [3]), .B(\array[113] [3]), .C(r_addr[0]), 
         .Z(n13520)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4978_3_lut.init = 16'hcaca;
    LUT4 i6316_3_lut (.A(\array[178] [0]), .B(\array[179] [0]), .C(r_addr[0]), 
         .Z(n14858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6316_3_lut.init = 16'hcaca;
    LUT4 i6315_3_lut (.A(\array[176] [0]), .B(\array[177] [0]), .C(r_addr[0]), 
         .Z(n14857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6315_3_lut.init = 16'hcaca;
    LUT4 i4977_3_lut (.A(\array[110] [3]), .B(\array[111] [3]), .C(r_addr[0]), 
         .Z(n13519)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4977_3_lut.init = 16'hcaca;
    LUT4 i4976_3_lut (.A(\array[108] [3]), .B(\array[109] [3]), .C(r_addr[0]), 
         .Z(n13518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4976_3_lut.init = 16'hcaca;
    LUT4 i4975_3_lut (.A(\array[106] [3]), .B(\array[107] [3]), .C(r_addr[0]), 
         .Z(n13517)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4975_3_lut.init = 16'hcaca;
    LUT4 i4974_3_lut (.A(\array[104] [3]), .B(\array[105] [3]), .C(r_addr[0]), 
         .Z(n13516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4974_3_lut.init = 16'hcaca;
    LUT4 i4973_3_lut (.A(\array[102] [3]), .B(\array[103] [3]), .C(r_addr[0]), 
         .Z(n13515)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4973_3_lut.init = 16'hcaca;
    LUT4 i4972_3_lut (.A(\array[100] [3]), .B(\array[101] [3]), .C(r_addr[0]), 
         .Z(n13514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4972_3_lut.init = 16'hcaca;
    LUT4 i4971_3_lut (.A(\array[98] [3]), .B(\array[99] [3]), .C(r_addr[0]), 
         .Z(n13513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4971_3_lut.init = 16'hcaca;
    LUT4 i4970_3_lut (.A(\array[96] [3]), .B(\array[97] [3]), .C(r_addr[0]), 
         .Z(n13512)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4970_3_lut.init = 16'hcaca;
    LUT4 i6229_3_lut (.A(\array[94] [0]), .B(\array[95] [0]), .C(r_addr[0]), 
         .Z(n14771)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6229_3_lut.init = 16'hcaca;
    LUT4 i6228_3_lut (.A(\array[92] [0]), .B(\array[93] [0]), .C(r_addr[0]), 
         .Z(n14770)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6228_3_lut.init = 16'hcaca;
    LUT4 i6227_3_lut (.A(\array[90] [0]), .B(\array[91] [0]), .C(r_addr[0]), 
         .Z(n14769)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6227_3_lut.init = 16'hcaca;
    LUT4 i6226_3_lut (.A(\array[88] [0]), .B(\array[89] [0]), .C(r_addr[0]), 
         .Z(n14768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6226_3_lut.init = 16'hcaca;
    LUT4 i6314_3_lut (.A(\array[174] [0]), .B(\array[175] [0]), .C(r_addr[0]), 
         .Z(n14856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6314_3_lut.init = 16'hcaca;
    LUT4 i6313_3_lut (.A(\array[172] [0]), .B(\array[173] [0]), .C(r_addr[0]), 
         .Z(n14855)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6313_3_lut.init = 16'hcaca;
    LUT4 i5688_3_lut (.A(\array[62] [6]), .B(\array[63] [6]), .C(r_addr[0]), 
         .Z(n14230)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5688_3_lut.init = 16'hcaca;
    LUT4 i5687_3_lut (.A(\array[60] [6]), .B(\array[61] [6]), .C(r_addr[0]), 
         .Z(n14229)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5687_3_lut.init = 16'hcaca;
    LUT4 i5686_3_lut (.A(\array[58] [6]), .B(\array[59] [6]), .C(r_addr[0]), 
         .Z(n14228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5686_3_lut.init = 16'hcaca;
    LUT4 i5685_3_lut (.A(\array[56] [6]), .B(\array[57] [6]), .C(r_addr[0]), 
         .Z(n14227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5685_3_lut.init = 16'hcaca;
    LUT4 i5684_3_lut (.A(\array[54] [6]), .B(\array[55] [6]), .C(r_addr[0]), 
         .Z(n14226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5684_3_lut.init = 16'hcaca;
    LUT4 i5683_3_lut (.A(\array[52] [6]), .B(\array[53] [6]), .C(r_addr[0]), 
         .Z(n14225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5683_3_lut.init = 16'hcaca;
    LUT4 i5682_3_lut (.A(\array[50] [6]), .B(\array[51] [6]), .C(r_addr[0]), 
         .Z(n14224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5682_3_lut.init = 16'hcaca;
    LUT4 i5681_3_lut (.A(\array[48] [6]), .B(\array[49] [6]), .C(r_addr[0]), 
         .Z(n14223)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5681_3_lut.init = 16'hcaca;
    LUT4 i6225_3_lut (.A(\array[86] [0]), .B(\array[87] [0]), .C(r_addr[0]), 
         .Z(n14767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6225_3_lut.init = 16'hcaca;
    LUT4 i6224_3_lut (.A(\array[84] [0]), .B(\array[85] [0]), .C(r_addr[0]), 
         .Z(n14766)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6224_3_lut.init = 16'hcaca;
    LUT4 i5680_3_lut (.A(\array[46] [6]), .B(\array[47] [6]), .C(r_addr[0]), 
         .Z(n14222)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5680_3_lut.init = 16'hcaca;
    LUT4 i5679_3_lut (.A(\array[44] [6]), .B(\array[45] [6]), .C(r_addr[0]), 
         .Z(n14221)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5679_3_lut.init = 16'hcaca;
    LUT4 i4954_3_lut (.A(\array[94] [3]), .B(\array[95] [3]), .C(r_addr[0]), 
         .Z(n13496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4954_3_lut.init = 16'hcaca;
    LUT4 i4953_3_lut (.A(\array[92] [3]), .B(\array[93] [3]), .C(r_addr[0]), 
         .Z(n13495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4953_3_lut.init = 16'hcaca;
    LUT4 i4952_3_lut (.A(\array[90] [3]), .B(\array[91] [3]), .C(r_addr[0]), 
         .Z(n13494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4952_3_lut.init = 16'hcaca;
    LUT4 i4951_3_lut (.A(\array[88] [3]), .B(\array[89] [3]), .C(r_addr[0]), 
         .Z(n13493)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4951_3_lut.init = 16'hcaca;
    LUT4 i5678_3_lut (.A(\array[42] [6]), .B(\array[43] [6]), .C(r_addr[0]), 
         .Z(n14220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5678_3_lut.init = 16'hcaca;
    LUT4 i5677_3_lut (.A(\array[40] [6]), .B(\array[41] [6]), .C(r_addr[0]), 
         .Z(n14219)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5677_3_lut.init = 16'hcaca;
    LUT4 i4950_3_lut (.A(\array[86] [3]), .B(\array[87] [3]), .C(r_addr[0]), 
         .Z(n13492)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4950_3_lut.init = 16'hcaca;
    LUT4 i4949_3_lut (.A(\array[84] [3]), .B(\array[85] [3]), .C(r_addr[0]), 
         .Z(n13491)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4949_3_lut.init = 16'hcaca;
    LUT4 i4948_3_lut (.A(\array[82] [3]), .B(\array[83] [3]), .C(r_addr[0]), 
         .Z(n13490)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4948_3_lut.init = 16'hcaca;
    LUT4 i4947_3_lut (.A(\array[80] [3]), .B(\array[81] [3]), .C(r_addr[0]), 
         .Z(n13489)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4947_3_lut.init = 16'hcaca;
    LUT4 i5676_3_lut (.A(\array[38] [6]), .B(\array[39] [6]), .C(r_addr[0]), 
         .Z(n14218)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5676_3_lut.init = 16'hcaca;
    LUT4 i5675_3_lut (.A(\array[36] [6]), .B(\array[37] [6]), .C(r_addr[0]), 
         .Z(n14217)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5675_3_lut.init = 16'hcaca;
    LUT4 i4946_3_lut (.A(\array[78] [3]), .B(\array[79] [3]), .C(r_addr[0]), 
         .Z(n13488)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4946_3_lut.init = 16'hcaca;
    LUT4 i4945_3_lut (.A(\array[76] [3]), .B(\array[77] [3]), .C(r_addr[0]), 
         .Z(n13487)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4945_3_lut.init = 16'hcaca;
    LUT4 i4944_3_lut (.A(\array[74] [3]), .B(\array[75] [3]), .C(r_addr[0]), 
         .Z(n13486)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4944_3_lut.init = 16'hcaca;
    LUT4 i4943_3_lut (.A(\array[72] [3]), .B(\array[73] [3]), .C(r_addr[0]), 
         .Z(n13485)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4943_3_lut.init = 16'hcaca;
    LUT4 i5674_3_lut (.A(\array[34] [6]), .B(\array[35] [6]), .C(r_addr[0]), 
         .Z(n14216)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5674_3_lut.init = 16'hcaca;
    LUT4 i5673_3_lut (.A(\array[32] [6]), .B(\array[33] [6]), .C(r_addr[0]), 
         .Z(n14215)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5673_3_lut.init = 16'hcaca;
    LUT4 i6223_3_lut (.A(\array[82] [0]), .B(\array[83] [0]), .C(r_addr[0]), 
         .Z(n14765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6223_3_lut.init = 16'hcaca;
    LUT4 i6222_3_lut (.A(\array[80] [0]), .B(\array[81] [0]), .C(r_addr[0]), 
         .Z(n14764)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6222_3_lut.init = 16'hcaca;
    LUT4 i6312_3_lut (.A(\array[170] [0]), .B(\array[171] [0]), .C(r_addr[0]), 
         .Z(n14854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6312_3_lut.init = 16'hcaca;
    LUT4 i6311_3_lut (.A(\array[168] [0]), .B(\array[169] [0]), .C(r_addr[0]), 
         .Z(n14853)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6311_3_lut.init = 16'hcaca;
    LUT4 i4942_3_lut (.A(\array[70] [3]), .B(\array[71] [3]), .C(r_addr[0]), 
         .Z(n13484)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4942_3_lut.init = 16'hcaca;
    LUT4 i4941_3_lut (.A(\array[68] [3]), .B(\array[69] [3]), .C(r_addr[0]), 
         .Z(n13483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4941_3_lut.init = 16'hcaca;
    LUT4 i4940_3_lut (.A(\array[66] [3]), .B(\array[67] [3]), .C(r_addr[0]), 
         .Z(n13482)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4940_3_lut.init = 16'hcaca;
    LUT4 i4939_3_lut (.A(\array[64] [3]), .B(\array[65] [3]), .C(r_addr[0]), 
         .Z(n13481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4939_3_lut.init = 16'hcaca;
    LUT4 i6221_3_lut (.A(\array[78] [0]), .B(\array[79] [0]), .C(r_addr[0]), 
         .Z(n14763)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6221_3_lut.init = 16'hcaca;
    LUT4 i6220_3_lut (.A(\array[76] [0]), .B(\array[77] [0]), .C(r_addr[0]), 
         .Z(n14762)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6220_3_lut.init = 16'hcaca;
    LUT4 i6219_3_lut (.A(\array[74] [0]), .B(\array[75] [0]), .C(r_addr[0]), 
         .Z(n14761)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6219_3_lut.init = 16'hcaca;
    LUT4 i6218_3_lut (.A(\array[72] [0]), .B(\array[73] [0]), .C(r_addr[0]), 
         .Z(n14760)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6218_3_lut.init = 16'hcaca;
    LUT4 i6310_3_lut (.A(\array[166] [0]), .B(\array[167] [0]), .C(r_addr[0]), 
         .Z(n14852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6310_3_lut.init = 16'hcaca;
    LUT4 i6309_3_lut (.A(\array[164] [0]), .B(\array[165] [0]), .C(r_addr[0]), 
         .Z(n14851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6309_3_lut.init = 16'hcaca;
    LUT4 i6217_3_lut (.A(\array[70] [0]), .B(\array[71] [0]), .C(r_addr[0]), 
         .Z(n14759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6217_3_lut.init = 16'hcaca;
    LUT4 i6216_3_lut (.A(\array[68] [0]), .B(\array[69] [0]), .C(r_addr[0]), 
         .Z(n14758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6216_3_lut.init = 16'hcaca;
    LUT4 i4923_3_lut (.A(\array[62] [3]), .B(\array[63] [3]), .C(r_addr[0]), 
         .Z(n13465)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4923_3_lut.init = 16'hcaca;
    LUT4 i4922_3_lut (.A(\array[60] [3]), .B(\array[61] [3]), .C(r_addr[0]), 
         .Z(n13464)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4922_3_lut.init = 16'hcaca;
    LUT4 i4921_3_lut (.A(\array[58] [3]), .B(\array[59] [3]), .C(r_addr[0]), 
         .Z(n13463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4921_3_lut.init = 16'hcaca;
    LUT4 i4920_3_lut (.A(\array[56] [3]), .B(\array[57] [3]), .C(r_addr[0]), 
         .Z(n13462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4920_3_lut.init = 16'hcaca;
    LUT4 i4919_3_lut (.A(\array[54] [3]), .B(\array[55] [3]), .C(r_addr[0]), 
         .Z(n13461)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4919_3_lut.init = 16'hcaca;
    LUT4 i4918_3_lut (.A(\array[52] [3]), .B(\array[53] [3]), .C(r_addr[0]), 
         .Z(n13460)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4918_3_lut.init = 16'hcaca;
    LUT4 i4917_3_lut (.A(\array[50] [3]), .B(\array[51] [3]), .C(r_addr[0]), 
         .Z(n13459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4917_3_lut.init = 16'hcaca;
    LUT4 i4916_3_lut (.A(\array[48] [3]), .B(\array[49] [3]), .C(r_addr[0]), 
         .Z(n13458)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4916_3_lut.init = 16'hcaca;
    LUT4 i4915_3_lut (.A(\array[46] [3]), .B(\array[47] [3]), .C(r_addr[0]), 
         .Z(n13457)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4915_3_lut.init = 16'hcaca;
    LUT4 i4914_3_lut (.A(\array[44] [3]), .B(\array[45] [3]), .C(r_addr[0]), 
         .Z(n13456)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4914_3_lut.init = 16'hcaca;
    LUT4 i4913_3_lut (.A(\array[42] [3]), .B(\array[43] [3]), .C(r_addr[0]), 
         .Z(n13455)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4913_3_lut.init = 16'hcaca;
    LUT4 i4912_3_lut (.A(\array[40] [3]), .B(\array[41] [3]), .C(r_addr[0]), 
         .Z(n13454)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4912_3_lut.init = 16'hcaca;
    LUT4 i4911_3_lut (.A(\array[38] [3]), .B(\array[39] [3]), .C(r_addr[0]), 
         .Z(n13453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4911_3_lut.init = 16'hcaca;
    LUT4 i4910_3_lut (.A(\array[36] [3]), .B(\array[37] [3]), .C(r_addr[0]), 
         .Z(n13452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4910_3_lut.init = 16'hcaca;
    LUT4 i6036_3_lut (.A(\array[158] [7]), .B(\array[159] [7]), .C(r_addr[0]), 
         .Z(n14578)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6036_3_lut.init = 16'hcaca;
    LUT4 i6035_3_lut (.A(\array[156] [7]), .B(\array[157] [7]), .C(r_addr[0]), 
         .Z(n14577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6035_3_lut.init = 16'hcaca;
    OB d_out_pad_7 (.I(d_out_c_7), .O(d_out[7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(21[26:31])
    LUT4 i6215_3_lut (.A(\array[66] [0]), .B(\array[67] [0]), .C(r_addr[0]), 
         .Z(n14757)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6215_3_lut.init = 16'hcaca;
    LUT4 i6214_3_lut (.A(\array[64] [0]), .B(\array[65] [0]), .C(r_addr[0]), 
         .Z(n14756)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6214_3_lut.init = 16'hcaca;
    VLO i7360 (.Z(GND_net));
    LUT4 i6308_3_lut (.A(\array[162] [0]), .B(\array[163] [0]), .C(r_addr[0]), 
         .Z(n14850)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6308_3_lut.init = 16'hcaca;
    LUT4 i6307_3_lut (.A(\array[160] [0]), .B(\array[161] [0]), .C(r_addr[0]), 
         .Z(n14849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6307_3_lut.init = 16'hcaca;
    LUT4 i4909_3_lut (.A(\array[34] [3]), .B(\array[35] [3]), .C(r_addr[0]), 
         .Z(n13451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4909_3_lut.init = 16'hcaca;
    LUT4 i4908_3_lut (.A(\array[32] [3]), .B(\array[33] [3]), .C(r_addr[0]), 
         .Z(n13450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4908_3_lut.init = 16'hcaca;
    LUT4 i6034_3_lut (.A(\array[154] [7]), .B(\array[155] [7]), .C(r_addr[0]), 
         .Z(n14576)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6034_3_lut.init = 16'hcaca;
    LUT4 i6033_3_lut (.A(\array[152] [7]), .B(\array[153] [7]), .C(r_addr[0]), 
         .Z(n14575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6033_3_lut.init = 16'hcaca;
    LUT4 i6032_3_lut (.A(\array[150] [7]), .B(\array[151] [7]), .C(r_addr[0]), 
         .Z(n14574)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6032_3_lut.init = 16'hcaca;
    LUT4 i6031_3_lut (.A(\array[148] [7]), .B(\array[149] [7]), .C(r_addr[0]), 
         .Z(n14573)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6031_3_lut.init = 16'hcaca;
    LUT4 i6030_3_lut (.A(\array[146] [7]), .B(\array[147] [7]), .C(r_addr[0]), 
         .Z(n14572)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6030_3_lut.init = 16'hcaca;
    LUT4 i6029_3_lut (.A(\array[144] [7]), .B(\array[145] [7]), .C(r_addr[0]), 
         .Z(n14571)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6029_3_lut.init = 16'hcaca;
    LUT4 i5657_3_lut (.A(\array[30] [6]), .B(\array[31] [6]), .C(r_addr[0]), 
         .Z(n14199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5657_3_lut.init = 16'hcaca;
    LUT4 i5656_3_lut (.A(\array[28] [6]), .B(\array[29] [6]), .C(r_addr[0]), 
         .Z(n14198)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5656_3_lut.init = 16'hcaca;
    LUT4 i5655_3_lut (.A(\array[26] [6]), .B(\array[27] [6]), .C(r_addr[0]), 
         .Z(n14197)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5655_3_lut.init = 16'hcaca;
    LUT4 i5654_3_lut (.A(\array[24] [6]), .B(\array[25] [6]), .C(r_addr[0]), 
         .Z(n14196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5654_3_lut.init = 16'hcaca;
    LUT4 i6028_3_lut (.A(\array[142] [7]), .B(\array[143] [7]), .C(r_addr[0]), 
         .Z(n14570)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6028_3_lut.init = 16'hcaca;
    LUT4 i6027_3_lut (.A(\array[140] [7]), .B(\array[141] [7]), .C(r_addr[0]), 
         .Z(n14569)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6027_3_lut.init = 16'hcaca;
    LUT4 i5653_3_lut (.A(\array[22] [6]), .B(\array[23] [6]), .C(r_addr[0]), 
         .Z(n14195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5653_3_lut.init = 16'hcaca;
    LUT4 i5652_3_lut (.A(\array[20] [6]), .B(\array[21] [6]), .C(r_addr[0]), 
         .Z(n14194)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5652_3_lut.init = 16'hcaca;
    LUT4 i5651_3_lut (.A(\array[18] [6]), .B(\array[19] [6]), .C(r_addr[0]), 
         .Z(n14193)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5651_3_lut.init = 16'hcaca;
    LUT4 i5650_3_lut (.A(\array[16] [6]), .B(\array[17] [6]), .C(r_addr[0]), 
         .Z(n14192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5650_3_lut.init = 16'hcaca;
    LUT4 i6026_3_lut (.A(\array[138] [7]), .B(\array[139] [7]), .C(r_addr[0]), 
         .Z(n14568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6026_3_lut.init = 16'hcaca;
    LUT4 i6025_3_lut (.A(\array[136] [7]), .B(\array[137] [7]), .C(r_addr[0]), 
         .Z(n14567)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6025_3_lut.init = 16'hcaca;
    LUT4 i5649_3_lut (.A(\array[14] [6]), .B(\array[15] [6]), .C(r_addr[0]), 
         .Z(n14191)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5649_3_lut.init = 16'hcaca;
    LUT4 i5648_3_lut (.A(\array[12] [6]), .B(\array[13] [6]), .C(r_addr[0]), 
         .Z(n14190)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5648_3_lut.init = 16'hcaca;
    LUT4 i4892_3_lut (.A(\array[30] [3]), .B(\array[31] [3]), .C(r_addr[0]), 
         .Z(n13434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4892_3_lut.init = 16'hcaca;
    LUT4 i4891_3_lut (.A(\array[28] [3]), .B(\array[29] [3]), .C(r_addr[0]), 
         .Z(n13433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4891_3_lut.init = 16'hcaca;
    LUT4 i5647_3_lut (.A(\array[10] [6]), .B(\array[11] [6]), .C(r_addr[0]), 
         .Z(n14189)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5647_3_lut.init = 16'hcaca;
    LUT4 i5646_3_lut (.A(\array[8] [6]), .B(\array[9] [6]), .C(r_addr[0]), 
         .Z(n14188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5646_3_lut.init = 16'hcaca;
    LUT4 i6024_3_lut (.A(\array[134] [7]), .B(\array[135] [7]), .C(r_addr[0]), 
         .Z(n14566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6024_3_lut.init = 16'hcaca;
    LUT4 i6023_3_lut (.A(\array[132] [7]), .B(\array[133] [7]), .C(r_addr[0]), 
         .Z(n14565)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6023_3_lut.init = 16'hcaca;
    LUT4 i4890_3_lut (.A(\array[26] [3]), .B(\array[27] [3]), .C(r_addr[0]), 
         .Z(n13432)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4890_3_lut.init = 16'hcaca;
    LUT4 i4889_3_lut (.A(\array[24] [3]), .B(\array[25] [3]), .C(r_addr[0]), 
         .Z(n13431)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4889_3_lut.init = 16'hcaca;
    LUT4 i4888_3_lut (.A(\array[22] [3]), .B(\array[23] [3]), .C(r_addr[0]), 
         .Z(n13430)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4888_3_lut.init = 16'hcaca;
    LUT4 i4887_3_lut (.A(\array[20] [3]), .B(\array[21] [3]), .C(r_addr[0]), 
         .Z(n13429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4887_3_lut.init = 16'hcaca;
    LUT4 i5645_3_lut (.A(\array[6] [6]), .B(\array[7] [6]), .C(r_addr[0]), 
         .Z(n14187)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5645_3_lut.init = 16'hcaca;
    LUT4 i5644_3_lut (.A(\array[4] [6]), .B(\array[5] [6]), .C(r_addr[0]), 
         .Z(n14186)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5644_3_lut.init = 16'hcaca;
    LUT4 i4886_3_lut (.A(\array[18] [3]), .B(\array[19] [3]), .C(r_addr[0]), 
         .Z(n13428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4886_3_lut.init = 16'hcaca;
    LUT4 i4885_3_lut (.A(\array[16] [3]), .B(\array[17] [3]), .C(r_addr[0]), 
         .Z(n13427)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4885_3_lut.init = 16'hcaca;
    LUT4 i4884_3_lut (.A(\array[14] [3]), .B(\array[15] [3]), .C(r_addr[0]), 
         .Z(n13426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4884_3_lut.init = 16'hcaca;
    LUT4 i4883_3_lut (.A(\array[12] [3]), .B(\array[13] [3]), .C(r_addr[0]), 
         .Z(n13425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4883_3_lut.init = 16'hcaca;
    LUT4 i5643_3_lut (.A(\array[2] [6]), .B(\array[3] [6]), .C(r_addr[0]), 
         .Z(n14185)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5643_3_lut.init = 16'hcaca;
    LUT4 i5642_3_lut (.A(\array[0] [6]), .B(\array[1] [6]), .C(r_addr[0]), 
         .Z(n14184)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5642_3_lut.init = 16'hcaca;
    LUT4 i6022_3_lut (.A(\array[130] [7]), .B(\array[131] [7]), .C(r_addr[0]), 
         .Z(n14564)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6022_3_lut.init = 16'hcaca;
    LUT4 i6021_3_lut (.A(\array[128] [7]), .B(\array[129] [7]), .C(r_addr[0]), 
         .Z(n14563)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6021_3_lut.init = 16'hcaca;
    LUT4 i4882_3_lut (.A(\array[10] [3]), .B(\array[11] [3]), .C(r_addr[0]), 
         .Z(n13424)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4882_3_lut.init = 16'hcaca;
    LUT4 i4881_3_lut (.A(\array[8] [3]), .B(\array[9] [3]), .C(r_addr[0]), 
         .Z(n13423)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4881_3_lut.init = 16'hcaca;
    LUT4 i4880_3_lut (.A(\array[6] [3]), .B(\array[7] [3]), .C(r_addr[0]), 
         .Z(n13422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4880_3_lut.init = 16'hcaca;
    LUT4 i4879_3_lut (.A(\array[4] [3]), .B(\array[5] [3]), .C(r_addr[0]), 
         .Z(n13421)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4879_3_lut.init = 16'hcaca;
    LUT4 i4878_3_lut (.A(\array[2] [3]), .B(\array[3] [3]), .C(r_addr[0]), 
         .Z(n13420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4878_3_lut.init = 16'hcaca;
    LUT4 i4877_3_lut (.A(\array[0] [3]), .B(\array[1] [3]), .C(r_addr[0]), 
         .Z(n13419)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4877_3_lut.init = 16'hcaca;
    LUT4 i6384_3_lut (.A(\array[254] [0]), .B(\array[255] [0]), .C(r_addr[0]), 
         .Z(n14926)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6384_3_lut.init = 16'hcaca;
    LUT4 i6383_3_lut (.A(\array[252] [0]), .B(\array[253] [0]), .C(r_addr[0]), 
         .Z(n14925)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6383_3_lut.init = 16'hcaca;
    LUT4 i4854_3_lut (.A(\array[254] [2]), .B(\array[255] [2]), .C(r_addr[0]), 
         .Z(n13396)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4854_3_lut.init = 16'hcaca;
    LUT4 i4853_3_lut (.A(\array[252] [2]), .B(\array[253] [2]), .C(r_addr[0]), 
         .Z(n13395)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4853_3_lut.init = 16'hcaca;
    LUT4 i4852_3_lut (.A(\array[250] [2]), .B(\array[251] [2]), .C(r_addr[0]), 
         .Z(n13394)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4852_3_lut.init = 16'hcaca;
    LUT4 i4851_3_lut (.A(\array[248] [2]), .B(\array[249] [2]), .C(r_addr[0]), 
         .Z(n13393)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4851_3_lut.init = 16'hcaca;
    LUT4 i4850_3_lut (.A(\array[246] [2]), .B(\array[247] [2]), .C(r_addr[0]), 
         .Z(n13392)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4850_3_lut.init = 16'hcaca;
    LUT4 i4849_3_lut (.A(\array[244] [2]), .B(\array[245] [2]), .C(r_addr[0]), 
         .Z(n13391)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4849_3_lut.init = 16'hcaca;
    LUT4 i4848_3_lut (.A(\array[242] [2]), .B(\array[243] [2]), .C(r_addr[0]), 
         .Z(n13390)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4848_3_lut.init = 16'hcaca;
    LUT4 i4847_3_lut (.A(\array[240] [2]), .B(\array[241] [2]), .C(r_addr[0]), 
         .Z(n13389)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4847_3_lut.init = 16'hcaca;
    LUT4 i4846_3_lut (.A(\array[238] [2]), .B(\array[239] [2]), .C(r_addr[0]), 
         .Z(n13388)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4846_3_lut.init = 16'hcaca;
    LUT4 i4845_3_lut (.A(\array[236] [2]), .B(\array[237] [2]), .C(r_addr[0]), 
         .Z(n13387)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4845_3_lut.init = 16'hcaca;
    LUT4 i4844_3_lut (.A(\array[234] [2]), .B(\array[235] [2]), .C(r_addr[0]), 
         .Z(n13386)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4844_3_lut.init = 16'hcaca;
    LUT4 i4843_3_lut (.A(\array[232] [2]), .B(\array[233] [2]), .C(r_addr[0]), 
         .Z(n13385)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4843_3_lut.init = 16'hcaca;
    LUT4 i4842_3_lut (.A(\array[230] [2]), .B(\array[231] [2]), .C(r_addr[0]), 
         .Z(n13384)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4842_3_lut.init = 16'hcaca;
    LUT4 i4841_3_lut (.A(\array[228] [2]), .B(\array[229] [2]), .C(r_addr[0]), 
         .Z(n13383)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4841_3_lut.init = 16'hcaca;
    LUT4 i4840_3_lut (.A(\array[226] [2]), .B(\array[227] [2]), .C(r_addr[0]), 
         .Z(n13382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4840_3_lut.init = 16'hcaca;
    LUT4 i4839_3_lut (.A(\array[224] [2]), .B(\array[225] [2]), .C(r_addr[0]), 
         .Z(n13381)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4839_3_lut.init = 16'hcaca;
    LUT4 i5619_3_lut (.A(\array[254] [5]), .B(\array[255] [5]), .C(r_addr[0]), 
         .Z(n14161)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5619_3_lut.init = 16'hcaca;
    LUT4 i5618_3_lut (.A(\array[252] [5]), .B(\array[253] [5]), .C(r_addr[0]), 
         .Z(n14160)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5618_3_lut.init = 16'hcaca;
    LUT4 i5617_3_lut (.A(\array[250] [5]), .B(\array[251] [5]), .C(r_addr[0]), 
         .Z(n14159)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5617_3_lut.init = 16'hcaca;
    LUT4 i5616_3_lut (.A(\array[248] [5]), .B(\array[249] [5]), .C(r_addr[0]), 
         .Z(n14158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5616_3_lut.init = 16'hcaca;
    LUT4 i4823_3_lut (.A(\array[222] [2]), .B(\array[223] [2]), .C(r_addr[0]), 
         .Z(n13365)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4823_3_lut.init = 16'hcaca;
    LUT4 i4822_3_lut (.A(\array[220] [2]), .B(\array[221] [2]), .C(r_addr[0]), 
         .Z(n13364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4822_3_lut.init = 16'hcaca;
    LUT4 i4821_3_lut (.A(\array[218] [2]), .B(\array[219] [2]), .C(r_addr[0]), 
         .Z(n13363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4821_3_lut.init = 16'hcaca;
    LUT4 i4820_3_lut (.A(\array[216] [2]), .B(\array[217] [2]), .C(r_addr[0]), 
         .Z(n13362)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4820_3_lut.init = 16'hcaca;
    LUT4 i5615_3_lut (.A(\array[246] [5]), .B(\array[247] [5]), .C(r_addr[0]), 
         .Z(n14157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5615_3_lut.init = 16'hcaca;
    LUT4 i5614_3_lut (.A(\array[244] [5]), .B(\array[245] [5]), .C(r_addr[0]), 
         .Z(n14156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5614_3_lut.init = 16'hcaca;
    LUT4 i4819_3_lut (.A(\array[214] [2]), .B(\array[215] [2]), .C(r_addr[0]), 
         .Z(n13361)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4819_3_lut.init = 16'hcaca;
    LUT4 i4818_3_lut (.A(\array[212] [2]), .B(\array[213] [2]), .C(r_addr[0]), 
         .Z(n13360)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4818_3_lut.init = 16'hcaca;
    LUT4 i4817_3_lut (.A(\array[210] [2]), .B(\array[211] [2]), .C(r_addr[0]), 
         .Z(n13359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4817_3_lut.init = 16'hcaca;
    LUT4 i4816_3_lut (.A(\array[208] [2]), .B(\array[209] [2]), .C(r_addr[0]), 
         .Z(n13358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4816_3_lut.init = 16'hcaca;
    LUT4 i5613_3_lut (.A(\array[242] [5]), .B(\array[243] [5]), .C(r_addr[0]), 
         .Z(n14155)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5613_3_lut.init = 16'hcaca;
    LUT4 i5612_3_lut (.A(\array[240] [5]), .B(\array[241] [5]), .C(r_addr[0]), 
         .Z(n14154)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5612_3_lut.init = 16'hcaca;
    LUT4 i4815_3_lut (.A(\array[206] [2]), .B(\array[207] [2]), .C(r_addr[0]), 
         .Z(n13357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4815_3_lut.init = 16'hcaca;
    LUT4 i4814_3_lut (.A(\array[204] [2]), .B(\array[205] [2]), .C(r_addr[0]), 
         .Z(n13356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4814_3_lut.init = 16'hcaca;
    LUT4 i4813_3_lut (.A(\array[202] [2]), .B(\array[203] [2]), .C(r_addr[0]), 
         .Z(n13355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4813_3_lut.init = 16'hcaca;
    LUT4 i4812_3_lut (.A(\array[200] [2]), .B(\array[201] [2]), .C(r_addr[0]), 
         .Z(n13354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4812_3_lut.init = 16'hcaca;
    LUT4 i5611_3_lut (.A(\array[238] [5]), .B(\array[239] [5]), .C(r_addr[0]), 
         .Z(n14153)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5611_3_lut.init = 16'hcaca;
    LUT4 i5610_3_lut (.A(\array[236] [5]), .B(\array[237] [5]), .C(r_addr[0]), 
         .Z(n14152)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5610_3_lut.init = 16'hcaca;
    LUT4 i6382_3_lut (.A(\array[250] [0]), .B(\array[251] [0]), .C(r_addr[0]), 
         .Z(n14924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6382_3_lut.init = 16'hcaca;
    LUT4 i6381_3_lut (.A(\array[248] [0]), .B(\array[249] [0]), .C(r_addr[0]), 
         .Z(n14923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6381_3_lut.init = 16'hcaca;
    LUT4 i4811_3_lut (.A(\array[198] [2]), .B(\array[199] [2]), .C(r_addr[0]), 
         .Z(n13353)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4811_3_lut.init = 16'hcaca;
    LUT4 i4810_3_lut (.A(\array[196] [2]), .B(\array[197] [2]), .C(r_addr[0]), 
         .Z(n13352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4810_3_lut.init = 16'hcaca;
    LUT4 i5609_3_lut (.A(\array[234] [5]), .B(\array[235] [5]), .C(r_addr[0]), 
         .Z(n14151)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5609_3_lut.init = 16'hcaca;
    LUT4 i5608_3_lut (.A(\array[232] [5]), .B(\array[233] [5]), .C(r_addr[0]), 
         .Z(n14150)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5608_3_lut.init = 16'hcaca;
    LUT4 i4809_3_lut (.A(\array[194] [2]), .B(\array[195] [2]), .C(r_addr[0]), 
         .Z(n13351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4809_3_lut.init = 16'hcaca;
    LUT4 i4808_3_lut (.A(\array[192] [2]), .B(\array[193] [2]), .C(r_addr[0]), 
         .Z(n13350)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4808_3_lut.init = 16'hcaca;
    LUT4 i5607_3_lut (.A(\array[230] [5]), .B(\array[231] [5]), .C(r_addr[0]), 
         .Z(n14149)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5607_3_lut.init = 16'hcaca;
    LUT4 i5606_3_lut (.A(\array[228] [5]), .B(\array[229] [5]), .C(r_addr[0]), 
         .Z(n14148)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5606_3_lut.init = 16'hcaca;
    LUT4 i5605_3_lut (.A(\array[226] [5]), .B(\array[227] [5]), .C(r_addr[0]), 
         .Z(n14147)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5605_3_lut.init = 16'hcaca;
    LUT4 i5604_3_lut (.A(\array[224] [5]), .B(\array[225] [5]), .C(r_addr[0]), 
         .Z(n14146)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5604_3_lut.init = 16'hcaca;
    LUT4 i6005_3_lut (.A(\array[126] [7]), .B(\array[127] [7]), .C(r_addr[0]), 
         .Z(n14547)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6005_3_lut.init = 16'hcaca;
    LUT4 i6004_3_lut (.A(\array[124] [7]), .B(\array[125] [7]), .C(r_addr[0]), 
         .Z(n14546)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6004_3_lut.init = 16'hcaca;
    LUT4 i4792_3_lut (.A(\array[190] [2]), .B(\array[191] [2]), .C(r_addr[0]), 
         .Z(n13334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4792_3_lut.init = 16'hcaca;
    LUT4 i4791_3_lut (.A(\array[188] [2]), .B(\array[189] [2]), .C(r_addr[0]), 
         .Z(n13333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4791_3_lut.init = 16'hcaca;
    IB addr_pad_0 (.I(addr[0]), .O(addr_c_0));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(19[27:31])
    IB addr_pad_1 (.I(addr[1]), .O(addr_c_1));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(19[27:31])
    IB addr_pad_2 (.I(addr[2]), .O(addr_c_2));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(19[27:31])
    IB addr_pad_3 (.I(addr[3]), .O(addr_c_3));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(19[27:31])
    IB addr_pad_4 (.I(addr[4]), .O(addr_c_4));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(19[27:31])
    IB addr_pad_5 (.I(addr[5]), .O(addr_c_5));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(19[27:31])
    IB addr_pad_6 (.I(addr[6]), .O(addr_c_6));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(19[27:31])
    IB addr_pad_7 (.I(addr[7]), .O(addr_c_7));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(19[27:31])
    IB d_in_pad_0 (.I(d_in[0]), .O(d_in_c_0));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(18[21:25])
    IB d_in_pad_1 (.I(d_in[1]), .O(d_in_c_1));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(18[21:25])
    IB d_in_pad_2 (.I(d_in[2]), .O(d_in_c_2));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(18[21:25])
    IB d_in_pad_3 (.I(d_in[3]), .O(d_in_c_3));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(18[21:25])
    IB d_in_pad_4 (.I(d_in[4]), .O(d_in_c_4));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(18[21:25])
    IB d_in_pad_5 (.I(d_in[5]), .O(d_in_c_5));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(18[21:25])
    IB d_in_pad_6 (.I(d_in[6]), .O(d_in_c_6));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(18[21:25])
    IB d_in_pad_7 (.I(d_in[7]), .O(d_in_c_7));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(18[21:25])
    IB clk_pad (.I(clk), .O(clk_c));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(17[30:33])
    IB rd_en_pad (.I(rd_en), .O(rd_en_c));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(17[23:28])
    IB wr_en_pad (.I(wr_en), .O(wr_en_c));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(17[16:21])
    OB d_out_pad_0 (.I(d_out_c_0), .O(d_out[0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(21[26:31])
    OB d_out_pad_1 (.I(d_out_c_1), .O(d_out[1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(21[26:31])
    OB d_out_pad_2 (.I(d_out_c_2), .O(d_out[2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(21[26:31])
    OB d_out_pad_3 (.I(d_out_c_3), .O(d_out[3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(21[26:31])
    OB d_out_pad_4 (.I(d_out_c_4), .O(d_out[4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(21[26:31])
    OB d_out_pad_5 (.I(d_out_c_5), .O(d_out[5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(21[26:31])
    OB d_out_pad_6 (.I(d_out_c_6), .O(d_out[6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(21[26:31])
    LUT4 i4790_3_lut (.A(\array[186] [2]), .B(\array[187] [2]), .C(r_addr[0]), 
         .Z(n13332)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4790_3_lut.init = 16'hcaca;
    LUT4 i4789_3_lut (.A(\array[184] [2]), .B(\array[185] [2]), .C(r_addr[0]), 
         .Z(n13331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4789_3_lut.init = 16'hcaca;
    LUT4 i4788_3_lut (.A(\array[182] [2]), .B(\array[183] [2]), .C(r_addr[0]), 
         .Z(n13330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4788_3_lut.init = 16'hcaca;
    LUT4 i4787_3_lut (.A(\array[180] [2]), .B(\array[181] [2]), .C(r_addr[0]), 
         .Z(n13329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4787_3_lut.init = 16'hcaca;
    LUT4 i6003_3_lut (.A(\array[122] [7]), .B(\array[123] [7]), .C(r_addr[0]), 
         .Z(n14545)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6003_3_lut.init = 16'hcaca;
    LUT4 i6002_3_lut (.A(\array[120] [7]), .B(\array[121] [7]), .C(r_addr[0]), 
         .Z(n14544)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6002_3_lut.init = 16'hcaca;
    FD1P3AX array_255___i1 (.D(array_0__7__N_4097[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[255] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1.GSR = "ENABLED";
    LUT4 mux_253_i4_3_lut_4_lut (.A(n15013), .B(n14992), .C(\array[6] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2105[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_253_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_253_i5_3_lut_4_lut (.A(n15013), .B(n14992), .C(\array[6] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2105[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_253_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_253_i6_3_lut_4_lut (.A(n15013), .B(n14992), .C(\array[6] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2105[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_253_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_253_i7_3_lut_4_lut (.A(n15013), .B(n14992), .C(\array[6] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2105[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_253_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_253_i8_3_lut_4_lut (.A(n15013), .B(n14992), .C(\array[6] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2105[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_253_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_252_i1_3_lut_4_lut (.A(n15014), .B(n14992), .C(\array[7] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2113[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_252_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_252_i2_3_lut_4_lut (.A(n15014), .B(n14992), .C(\array[7] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2113[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_252_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_220_i1_3_lut_4_lut (.A(n15014), .B(n14994), .C(\array[39] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2369[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_220_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5329_3_lut (.A(\array[214] [4]), .B(\array[215] [4]), .C(r_addr[0]), 
         .Z(n13871)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5329_3_lut.init = 16'hcaca;
    LUT4 i5328_3_lut (.A(\array[212] [4]), .B(\array[213] [4]), .C(r_addr[0]), 
         .Z(n13870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5328_3_lut.init = 16'hcaca;
    LUT4 i5872_3_lut (.A(\array[250] [6]), .B(\array[251] [6]), .C(r_addr[0]), 
         .Z(n14414)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5872_3_lut.init = 16'hcaca;
    LUT4 i5871_3_lut (.A(\array[248] [6]), .B(\array[249] [6]), .C(r_addr[0]), 
         .Z(n14413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5871_3_lut.init = 16'hcaca;
    LUT4 i5327_3_lut (.A(\array[210] [4]), .B(\array[211] [4]), .C(r_addr[0]), 
         .Z(n13869)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5327_3_lut.init = 16'hcaca;
    LUT4 i5326_3_lut (.A(\array[208] [4]), .B(\array[209] [4]), .C(r_addr[0]), 
         .Z(n13868)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5326_3_lut.init = 16'hcaca;
    LUT4 i5325_3_lut (.A(\array[206] [4]), .B(\array[207] [4]), .C(r_addr[0]), 
         .Z(n13867)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5325_3_lut.init = 16'hcaca;
    LUT4 i5324_3_lut (.A(\array[204] [4]), .B(\array[205] [4]), .C(r_addr[0]), 
         .Z(n13866)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5324_3_lut.init = 16'hcaca;
    LUT4 i5870_3_lut (.A(\array[246] [6]), .B(\array[247] [6]), .C(r_addr[0]), 
         .Z(n14412)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5870_3_lut.init = 16'hcaca;
    LUT4 i5869_3_lut (.A(\array[244] [6]), .B(\array[245] [6]), .C(r_addr[0]), 
         .Z(n14411)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5869_3_lut.init = 16'hcaca;
    LUT4 i5323_3_lut (.A(\array[202] [4]), .B(\array[203] [4]), .C(r_addr[0]), 
         .Z(n13865)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5323_3_lut.init = 16'hcaca;
    LUT4 i5322_3_lut (.A(\array[200] [4]), .B(\array[201] [4]), .C(r_addr[0]), 
         .Z(n13864)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5322_3_lut.init = 16'hcaca;
    LUT4 i5321_3_lut (.A(\array[198] [4]), .B(\array[199] [4]), .C(r_addr[0]), 
         .Z(n13863)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5321_3_lut.init = 16'hcaca;
    LUT4 i5320_3_lut (.A(\array[196] [4]), .B(\array[197] [4]), .C(r_addr[0]), 
         .Z(n13862)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5320_3_lut.init = 16'hcaca;
    LUT4 i5868_3_lut (.A(\array[242] [6]), .B(\array[243] [6]), .C(r_addr[0]), 
         .Z(n14410)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5868_3_lut.init = 16'hcaca;
    LUT4 i5867_3_lut (.A(\array[240] [6]), .B(\array[241] [6]), .C(r_addr[0]), 
         .Z(n14409)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5867_3_lut.init = 16'hcaca;
    LUT4 i5319_3_lut (.A(\array[194] [4]), .B(\array[195] [4]), .C(r_addr[0]), 
         .Z(n13861)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5319_3_lut.init = 16'hcaca;
    LUT4 i5318_3_lut (.A(\array[192] [4]), .B(\array[193] [4]), .C(r_addr[0]), 
         .Z(n13860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5318_3_lut.init = 16'hcaca;
    LUT4 i5866_3_lut (.A(\array[238] [6]), .B(\array[239] [6]), .C(r_addr[0]), 
         .Z(n14408)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5866_3_lut.init = 16'hcaca;
    LUT4 i5865_3_lut (.A(\array[236] [6]), .B(\array[237] [6]), .C(r_addr[0]), 
         .Z(n14407)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5865_3_lut.init = 16'hcaca;
    LUT4 i5864_3_lut (.A(\array[234] [6]), .B(\array[235] [6]), .C(r_addr[0]), 
         .Z(n14406)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5864_3_lut.init = 16'hcaca;
    LUT4 i5863_3_lut (.A(\array[232] [6]), .B(\array[233] [6]), .C(r_addr[0]), 
         .Z(n14405)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5863_3_lut.init = 16'hcaca;
    LUT4 i5862_3_lut (.A(\array[230] [6]), .B(\array[231] [6]), .C(r_addr[0]), 
         .Z(n14404)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5862_3_lut.init = 16'hcaca;
    LUT4 i5861_3_lut (.A(\array[228] [6]), .B(\array[229] [6]), .C(r_addr[0]), 
         .Z(n14403)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5861_3_lut.init = 16'hcaca;
    LUT4 i5860_3_lut (.A(\array[226] [6]), .B(\array[227] [6]), .C(r_addr[0]), 
         .Z(n14402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5860_3_lut.init = 16'hcaca;
    LUT4 i5859_3_lut (.A(\array[224] [6]), .B(\array[225] [6]), .C(r_addr[0]), 
         .Z(n14401)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5859_3_lut.init = 16'hcaca;
    LUT4 i5302_3_lut (.A(\array[190] [4]), .B(\array[191] [4]), .C(r_addr[0]), 
         .Z(n13844)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5302_3_lut.init = 16'hcaca;
    LUT4 i5301_3_lut (.A(\array[188] [4]), .B(\array[189] [4]), .C(r_addr[0]), 
         .Z(n13843)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5301_3_lut.init = 16'hcaca;
    LUT4 i5300_3_lut (.A(\array[186] [4]), .B(\array[187] [4]), .C(r_addr[0]), 
         .Z(n13842)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5300_3_lut.init = 16'hcaca;
    LUT4 i5299_3_lut (.A(\array[184] [4]), .B(\array[185] [4]), .C(r_addr[0]), 
         .Z(n13841)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5299_3_lut.init = 16'hcaca;
    LUT4 i5298_3_lut (.A(\array[182] [4]), .B(\array[183] [4]), .C(r_addr[0]), 
         .Z(n13840)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5298_3_lut.init = 16'hcaca;
    LUT4 i5297_3_lut (.A(\array[180] [4]), .B(\array[181] [4]), .C(r_addr[0]), 
         .Z(n13839)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5297_3_lut.init = 16'hcaca;
    LUT4 i5296_3_lut (.A(\array[178] [4]), .B(\array[179] [4]), .C(r_addr[0]), 
         .Z(n13838)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5296_3_lut.init = 16'hcaca;
    LUT4 i5295_3_lut (.A(\array[176] [4]), .B(\array[177] [4]), .C(r_addr[0]), 
         .Z(n13837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5295_3_lut.init = 16'hcaca;
    LUT4 i5294_3_lut (.A(\array[174] [4]), .B(\array[175] [4]), .C(r_addr[0]), 
         .Z(n13836)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5294_3_lut.init = 16'hcaca;
    LUT4 i5293_3_lut (.A(\array[172] [4]), .B(\array[173] [4]), .C(r_addr[0]), 
         .Z(n13835)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5293_3_lut.init = 16'hcaca;
    LUT4 i5292_3_lut (.A(\array[170] [4]), .B(\array[171] [4]), .C(r_addr[0]), 
         .Z(n13834)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5292_3_lut.init = 16'hcaca;
    LUT4 i5291_3_lut (.A(\array[168] [4]), .B(\array[169] [4]), .C(r_addr[0]), 
         .Z(n13833)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5291_3_lut.init = 16'hcaca;
    LUT4 i5290_3_lut (.A(\array[166] [4]), .B(\array[167] [4]), .C(r_addr[0]), 
         .Z(n13832)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5290_3_lut.init = 16'hcaca;
    LUT4 i5289_3_lut (.A(\array[164] [4]), .B(\array[165] [4]), .C(r_addr[0]), 
         .Z(n13831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5289_3_lut.init = 16'hcaca;
    LUT4 i5288_3_lut (.A(\array[162] [4]), .B(\array[163] [4]), .C(r_addr[0]), 
         .Z(n13830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5288_3_lut.init = 16'hcaca;
    LUT4 i5287_3_lut (.A(\array[160] [4]), .B(\array[161] [4]), .C(r_addr[0]), 
         .Z(n13829)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5287_3_lut.init = 16'hcaca;
    LUT4 i6129_3_lut (.A(\array[254] [7]), .B(\array[255] [7]), .C(r_addr[0]), 
         .Z(n14671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6129_3_lut.init = 16'hcaca;
    LUT4 i6128_3_lut (.A(\array[252] [7]), .B(\array[253] [7]), .C(r_addr[0]), 
         .Z(n14670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6128_3_lut.init = 16'hcaca;
    LUT4 i6127_3_lut (.A(\array[250] [7]), .B(\array[251] [7]), .C(r_addr[0]), 
         .Z(n14669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6127_3_lut.init = 16'hcaca;
    LUT4 i6126_3_lut (.A(\array[248] [7]), .B(\array[249] [7]), .C(r_addr[0]), 
         .Z(n14668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6126_3_lut.init = 16'hcaca;
    LUT4 i6125_3_lut (.A(\array[246] [7]), .B(\array[247] [7]), .C(r_addr[0]), 
         .Z(n14667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6125_3_lut.init = 16'hcaca;
    LUT4 i6124_3_lut (.A(\array[244] [7]), .B(\array[245] [7]), .C(r_addr[0]), 
         .Z(n14666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6124_3_lut.init = 16'hcaca;
    LUT4 i6123_3_lut (.A(\array[242] [7]), .B(\array[243] [7]), .C(r_addr[0]), 
         .Z(n14665)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6123_3_lut.init = 16'hcaca;
    LUT4 i6122_3_lut (.A(\array[240] [7]), .B(\array[241] [7]), .C(r_addr[0]), 
         .Z(n14664)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6122_3_lut.init = 16'hcaca;
    LUT4 i5271_3_lut (.A(\array[158] [4]), .B(\array[159] [4]), .C(r_addr[0]), 
         .Z(n13813)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5271_3_lut.init = 16'hcaca;
    LUT4 i5270_3_lut (.A(\array[156] [4]), .B(\array[157] [4]), .C(r_addr[0]), 
         .Z(n13812)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5270_3_lut.init = 16'hcaca;
    LUT4 i5843_3_lut (.A(\array[222] [6]), .B(\array[223] [6]), .C(r_addr[0]), 
         .Z(n14385)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5843_3_lut.init = 16'hcaca;
    LUT4 i5842_3_lut (.A(\array[220] [6]), .B(\array[221] [6]), .C(r_addr[0]), 
         .Z(n14384)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5842_3_lut.init = 16'hcaca;
    LUT4 i5269_3_lut (.A(\array[154] [4]), .B(\array[155] [4]), .C(r_addr[0]), 
         .Z(n13811)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5269_3_lut.init = 16'hcaca;
    LUT4 i5268_3_lut (.A(\array[152] [4]), .B(\array[153] [4]), .C(r_addr[0]), 
         .Z(n13810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5268_3_lut.init = 16'hcaca;
    LUT4 i5267_3_lut (.A(\array[150] [4]), .B(\array[151] [4]), .C(r_addr[0]), 
         .Z(n13809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5267_3_lut.init = 16'hcaca;
    LUT4 i5266_3_lut (.A(\array[148] [4]), .B(\array[149] [4]), .C(r_addr[0]), 
         .Z(n13808)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5266_3_lut.init = 16'hcaca;
    LUT4 i5841_3_lut (.A(\array[218] [6]), .B(\array[219] [6]), .C(r_addr[0]), 
         .Z(n14383)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5841_3_lut.init = 16'hcaca;
    LUT4 i5840_3_lut (.A(\array[216] [6]), .B(\array[217] [6]), .C(r_addr[0]), 
         .Z(n14382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5840_3_lut.init = 16'hcaca;
    LUT4 i6121_3_lut (.A(\array[238] [7]), .B(\array[239] [7]), .C(r_addr[0]), 
         .Z(n14663)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6121_3_lut.init = 16'hcaca;
    LUT4 i6120_3_lut (.A(\array[236] [7]), .B(\array[237] [7]), .C(r_addr[0]), 
         .Z(n14662)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6120_3_lut.init = 16'hcaca;
    LUT4 i5265_3_lut (.A(\array[146] [4]), .B(\array[147] [4]), .C(r_addr[0]), 
         .Z(n13807)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5265_3_lut.init = 16'hcaca;
    LUT4 i5264_3_lut (.A(\array[144] [4]), .B(\array[145] [4]), .C(r_addr[0]), 
         .Z(n13806)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5264_3_lut.init = 16'hcaca;
    LUT4 i5263_3_lut (.A(\array[142] [4]), .B(\array[143] [4]), .C(r_addr[0]), 
         .Z(n13805)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5263_3_lut.init = 16'hcaca;
    LUT4 i5262_3_lut (.A(\array[140] [4]), .B(\array[141] [4]), .C(r_addr[0]), 
         .Z(n13804)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5262_3_lut.init = 16'hcaca;
    LUT4 i5839_3_lut (.A(\array[214] [6]), .B(\array[215] [6]), .C(r_addr[0]), 
         .Z(n14381)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5839_3_lut.init = 16'hcaca;
    LUT4 i5838_3_lut (.A(\array[212] [6]), .B(\array[213] [6]), .C(r_addr[0]), 
         .Z(n14380)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5838_3_lut.init = 16'hcaca;
    LUT4 i5261_3_lut (.A(\array[138] [4]), .B(\array[139] [4]), .C(r_addr[0]), 
         .Z(n13803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5261_3_lut.init = 16'hcaca;
    LUT4 i5260_3_lut (.A(\array[136] [4]), .B(\array[137] [4]), .C(r_addr[0]), 
         .Z(n13802)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5260_3_lut.init = 16'hcaca;
    LUT4 i5259_3_lut (.A(\array[134] [4]), .B(\array[135] [4]), .C(r_addr[0]), 
         .Z(n13801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5259_3_lut.init = 16'hcaca;
    LUT4 i5258_3_lut (.A(\array[132] [4]), .B(\array[133] [4]), .C(r_addr[0]), 
         .Z(n13800)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5258_3_lut.init = 16'hcaca;
    LUT4 i5837_3_lut (.A(\array[210] [6]), .B(\array[211] [6]), .C(r_addr[0]), 
         .Z(n14379)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5837_3_lut.init = 16'hcaca;
    LUT4 i5836_3_lut (.A(\array[208] [6]), .B(\array[209] [6]), .C(r_addr[0]), 
         .Z(n14378)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5836_3_lut.init = 16'hcaca;
    LUT4 i6119_3_lut (.A(\array[234] [7]), .B(\array[235] [7]), .C(r_addr[0]), 
         .Z(n14661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6119_3_lut.init = 16'hcaca;
    LUT4 i6118_3_lut (.A(\array[232] [7]), .B(\array[233] [7]), .C(r_addr[0]), 
         .Z(n14660)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6118_3_lut.init = 16'hcaca;
    LUT4 i5257_3_lut (.A(\array[130] [4]), .B(\array[131] [4]), .C(r_addr[0]), 
         .Z(n13799)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5257_3_lut.init = 16'hcaca;
    LUT4 i5256_3_lut (.A(\array[128] [4]), .B(\array[129] [4]), .C(r_addr[0]), 
         .Z(n13798)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5256_3_lut.init = 16'hcaca;
    LUT4 i5835_3_lut (.A(\array[206] [6]), .B(\array[207] [6]), .C(r_addr[0]), 
         .Z(n14377)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5835_3_lut.init = 16'hcaca;
    LUT4 i5834_3_lut (.A(\array[204] [6]), .B(\array[205] [6]), .C(r_addr[0]), 
         .Z(n14376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5834_3_lut.init = 16'hcaca;
    LUT4 i5833_3_lut (.A(\array[202] [6]), .B(\array[203] [6]), .C(r_addr[0]), 
         .Z(n14375)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5833_3_lut.init = 16'hcaca;
    LUT4 i5832_3_lut (.A(\array[200] [6]), .B(\array[201] [6]), .C(r_addr[0]), 
         .Z(n14374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5832_3_lut.init = 16'hcaca;
    LUT4 i6117_3_lut (.A(\array[230] [7]), .B(\array[231] [7]), .C(r_addr[0]), 
         .Z(n14659)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6117_3_lut.init = 16'hcaca;
    LUT4 i6116_3_lut (.A(\array[228] [7]), .B(\array[229] [7]), .C(r_addr[0]), 
         .Z(n14658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6116_3_lut.init = 16'hcaca;
    LUT4 i5831_3_lut (.A(\array[198] [6]), .B(\array[199] [6]), .C(r_addr[0]), 
         .Z(n14373)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5831_3_lut.init = 16'hcaca;
    LUT4 i5830_3_lut (.A(\array[196] [6]), .B(\array[197] [6]), .C(r_addr[0]), 
         .Z(n14372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5830_3_lut.init = 16'hcaca;
    LUT4 i5829_3_lut (.A(\array[194] [6]), .B(\array[195] [6]), .C(r_addr[0]), 
         .Z(n14371)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5829_3_lut.init = 16'hcaca;
    LUT4 i5828_3_lut (.A(\array[192] [6]), .B(\array[193] [6]), .C(r_addr[0]), 
         .Z(n14370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5828_3_lut.init = 16'hcaca;
    LUT4 i6115_3_lut (.A(\array[226] [7]), .B(\array[227] [7]), .C(r_addr[0]), 
         .Z(n14657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6115_3_lut.init = 16'hcaca;
    LUT4 i6114_3_lut (.A(\array[224] [7]), .B(\array[225] [7]), .C(r_addr[0]), 
         .Z(n14656)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6114_3_lut.init = 16'hcaca;
    LUT4 i5240_3_lut (.A(\array[126] [4]), .B(\array[127] [4]), .C(r_addr[0]), 
         .Z(n13782)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5240_3_lut.init = 16'hcaca;
    LUT4 i5239_3_lut (.A(\array[124] [4]), .B(\array[125] [4]), .C(r_addr[0]), 
         .Z(n13781)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5239_3_lut.init = 16'hcaca;
    LUT4 i5238_3_lut (.A(\array[122] [4]), .B(\array[123] [4]), .C(r_addr[0]), 
         .Z(n13780)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5238_3_lut.init = 16'hcaca;
    LUT4 i5237_3_lut (.A(\array[120] [4]), .B(\array[121] [4]), .C(r_addr[0]), 
         .Z(n13779)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5237_3_lut.init = 16'hcaca;
    LUT4 i5236_3_lut (.A(\array[118] [4]), .B(\array[119] [4]), .C(r_addr[0]), 
         .Z(n13778)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5236_3_lut.init = 16'hcaca;
    LUT4 i5235_3_lut (.A(\array[116] [4]), .B(\array[117] [4]), .C(r_addr[0]), 
         .Z(n13777)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5235_3_lut.init = 16'hcaca;
    LUT4 i5234_3_lut (.A(\array[114] [4]), .B(\array[115] [4]), .C(r_addr[0]), 
         .Z(n13776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5234_3_lut.init = 16'hcaca;
    LUT4 i5233_3_lut (.A(\array[112] [4]), .B(\array[113] [4]), .C(r_addr[0]), 
         .Z(n13775)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5233_3_lut.init = 16'hcaca;
    LUT4 i5232_3_lut (.A(\array[110] [4]), .B(\array[111] [4]), .C(r_addr[0]), 
         .Z(n13774)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5232_3_lut.init = 16'hcaca;
    LUT4 i5231_3_lut (.A(\array[108] [4]), .B(\array[109] [4]), .C(r_addr[0]), 
         .Z(n13773)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5231_3_lut.init = 16'hcaca;
    LUT4 i5230_3_lut (.A(\array[106] [4]), .B(\array[107] [4]), .C(r_addr[0]), 
         .Z(n13772)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5230_3_lut.init = 16'hcaca;
    LUT4 i5229_3_lut (.A(\array[104] [4]), .B(\array[105] [4]), .C(r_addr[0]), 
         .Z(n13771)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5229_3_lut.init = 16'hcaca;
    LUT4 i5228_3_lut (.A(\array[102] [4]), .B(\array[103] [4]), .C(r_addr[0]), 
         .Z(n13770)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5228_3_lut.init = 16'hcaca;
    LUT4 i5227_3_lut (.A(\array[100] [4]), .B(\array[101] [4]), .C(r_addr[0]), 
         .Z(n13769)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5227_3_lut.init = 16'hcaca;
    LUT4 i5226_3_lut (.A(\array[98] [4]), .B(\array[99] [4]), .C(r_addr[0]), 
         .Z(n13768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5226_3_lut.init = 16'hcaca;
    LUT4 i5225_3_lut (.A(\array[96] [4]), .B(\array[97] [4]), .C(r_addr[0]), 
         .Z(n13767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5225_3_lut.init = 16'hcaca;
    LUT4 i6260_3_lut (.A(\array[126] [0]), .B(\array[127] [0]), .C(r_addr[0]), 
         .Z(n14802)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6260_3_lut.init = 16'hcaca;
    LUT4 i6259_3_lut (.A(\array[124] [0]), .B(\array[125] [0]), .C(r_addr[0]), 
         .Z(n14801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6259_3_lut.init = 16'hcaca;
    LUT4 i6258_3_lut (.A(\array[122] [0]), .B(\array[123] [0]), .C(r_addr[0]), 
         .Z(n14800)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6258_3_lut.init = 16'hcaca;
    LUT4 i6257_3_lut (.A(\array[120] [0]), .B(\array[121] [0]), .C(r_addr[0]), 
         .Z(n14799)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6257_3_lut.init = 16'hcaca;
    LUT4 i5812_3_lut (.A(\array[190] [6]), .B(\array[191] [6]), .C(r_addr[0]), 
         .Z(n14354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5812_3_lut.init = 16'hcaca;
    LUT4 i5811_3_lut (.A(\array[188] [6]), .B(\array[189] [6]), .C(r_addr[0]), 
         .Z(n14353)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5811_3_lut.init = 16'hcaca;
    LUT4 i5209_3_lut (.A(\array[94] [4]), .B(\array[95] [4]), .C(r_addr[0]), 
         .Z(n13751)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5209_3_lut.init = 16'hcaca;
    LUT4 i5208_3_lut (.A(\array[92] [4]), .B(\array[93] [4]), .C(r_addr[0]), 
         .Z(n13750)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5208_3_lut.init = 16'hcaca;
    LUT4 i5207_3_lut (.A(\array[90] [4]), .B(\array[91] [4]), .C(r_addr[0]), 
         .Z(n13749)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5207_3_lut.init = 16'hcaca;
    LUT4 i5206_3_lut (.A(\array[88] [4]), .B(\array[89] [4]), .C(r_addr[0]), 
         .Z(n13748)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5206_3_lut.init = 16'hcaca;
    LUT4 i5810_3_lut (.A(\array[186] [6]), .B(\array[187] [6]), .C(r_addr[0]), 
         .Z(n14352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5810_3_lut.init = 16'hcaca;
    LUT4 i5809_3_lut (.A(\array[184] [6]), .B(\array[185] [6]), .C(r_addr[0]), 
         .Z(n14351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5809_3_lut.init = 16'hcaca;
    LUT4 i5205_3_lut (.A(\array[86] [4]), .B(\array[87] [4]), .C(r_addr[0]), 
         .Z(n13747)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5205_3_lut.init = 16'hcaca;
    LUT4 i5204_3_lut (.A(\array[84] [4]), .B(\array[85] [4]), .C(r_addr[0]), 
         .Z(n13746)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5204_3_lut.init = 16'hcaca;
    LUT4 i5203_3_lut (.A(\array[82] [4]), .B(\array[83] [4]), .C(r_addr[0]), 
         .Z(n13745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5203_3_lut.init = 16'hcaca;
    LUT4 i5202_3_lut (.A(\array[80] [4]), .B(\array[81] [4]), .C(r_addr[0]), 
         .Z(n13744)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5202_3_lut.init = 16'hcaca;
    LUT4 i5808_3_lut (.A(\array[182] [6]), .B(\array[183] [6]), .C(r_addr[0]), 
         .Z(n14350)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5808_3_lut.init = 16'hcaca;
    LUT4 i5807_3_lut (.A(\array[180] [6]), .B(\array[181] [6]), .C(r_addr[0]), 
         .Z(n14349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5807_3_lut.init = 16'hcaca;
    LUT4 i5201_3_lut (.A(\array[78] [4]), .B(\array[79] [4]), .C(r_addr[0]), 
         .Z(n13743)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5201_3_lut.init = 16'hcaca;
    LUT4 i5200_3_lut (.A(\array[76] [4]), .B(\array[77] [4]), .C(r_addr[0]), 
         .Z(n13742)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5200_3_lut.init = 16'hcaca;
    LUT4 i5199_3_lut (.A(\array[74] [4]), .B(\array[75] [4]), .C(r_addr[0]), 
         .Z(n13741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5199_3_lut.init = 16'hcaca;
    LUT4 i5198_3_lut (.A(\array[72] [4]), .B(\array[73] [4]), .C(r_addr[0]), 
         .Z(n13740)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5198_3_lut.init = 16'hcaca;
    LUT4 i5806_3_lut (.A(\array[178] [6]), .B(\array[179] [6]), .C(r_addr[0]), 
         .Z(n14348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5806_3_lut.init = 16'hcaca;
    LUT4 i5805_3_lut (.A(\array[176] [6]), .B(\array[177] [6]), .C(r_addr[0]), 
         .Z(n14347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5805_3_lut.init = 16'hcaca;
    LUT4 i6256_3_lut (.A(\array[118] [0]), .B(\array[119] [0]), .C(r_addr[0]), 
         .Z(n14798)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6256_3_lut.init = 16'hcaca;
    LUT4 i6255_3_lut (.A(\array[116] [0]), .B(\array[117] [0]), .C(r_addr[0]), 
         .Z(n14797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6255_3_lut.init = 16'hcaca;
    LUT4 i5197_3_lut (.A(\array[70] [4]), .B(\array[71] [4]), .C(r_addr[0]), 
         .Z(n13739)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5197_3_lut.init = 16'hcaca;
    LUT4 i5196_3_lut (.A(\array[68] [4]), .B(\array[69] [4]), .C(r_addr[0]), 
         .Z(n13738)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5196_3_lut.init = 16'hcaca;
    LUT4 i5195_3_lut (.A(\array[66] [4]), .B(\array[67] [4]), .C(r_addr[0]), 
         .Z(n13737)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5195_3_lut.init = 16'hcaca;
    LUT4 i5194_3_lut (.A(\array[64] [4]), .B(\array[65] [4]), .C(r_addr[0]), 
         .Z(n13736)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5194_3_lut.init = 16'hcaca;
    LUT4 i5804_3_lut (.A(\array[174] [6]), .B(\array[175] [6]), .C(r_addr[0]), 
         .Z(n14346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5804_3_lut.init = 16'hcaca;
    LUT4 i5803_3_lut (.A(\array[172] [6]), .B(\array[173] [6]), .C(r_addr[0]), 
         .Z(n14345)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5803_3_lut.init = 16'hcaca;
    LUT4 i5802_3_lut (.A(\array[170] [6]), .B(\array[171] [6]), .C(r_addr[0]), 
         .Z(n14344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5802_3_lut.init = 16'hcaca;
    LUT4 i5801_3_lut (.A(\array[168] [6]), .B(\array[169] [6]), .C(r_addr[0]), 
         .Z(n14343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5801_3_lut.init = 16'hcaca;
    LUT4 i5800_3_lut (.A(\array[166] [6]), .B(\array[167] [6]), .C(r_addr[0]), 
         .Z(n14342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5800_3_lut.init = 16'hcaca;
    LUT4 i5799_3_lut (.A(\array[164] [6]), .B(\array[165] [6]), .C(r_addr[0]), 
         .Z(n14341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5799_3_lut.init = 16'hcaca;
    LUT4 i5798_3_lut (.A(\array[162] [6]), .B(\array[163] [6]), .C(r_addr[0]), 
         .Z(n14340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5798_3_lut.init = 16'hcaca;
    LUT4 i5797_3_lut (.A(\array[160] [6]), .B(\array[161] [6]), .C(r_addr[0]), 
         .Z(n14339)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5797_3_lut.init = 16'hcaca;
    LUT4 i6254_3_lut (.A(\array[114] [0]), .B(\array[115] [0]), .C(r_addr[0]), 
         .Z(n14796)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6254_3_lut.init = 16'hcaca;
    LUT4 i6253_3_lut (.A(\array[112] [0]), .B(\array[113] [0]), .C(r_addr[0]), 
         .Z(n14795)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6253_3_lut.init = 16'hcaca;
    LUT4 i6252_3_lut (.A(\array[110] [0]), .B(\array[111] [0]), .C(r_addr[0]), 
         .Z(n14794)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6252_3_lut.init = 16'hcaca;
    LUT4 i6251_3_lut (.A(\array[108] [0]), .B(\array[109] [0]), .C(r_addr[0]), 
         .Z(n14793)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6251_3_lut.init = 16'hcaca;
    LUT4 i6250_3_lut (.A(\array[106] [0]), .B(\array[107] [0]), .C(r_addr[0]), 
         .Z(n14792)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6250_3_lut.init = 16'hcaca;
    LUT4 i6249_3_lut (.A(\array[104] [0]), .B(\array[105] [0]), .C(r_addr[0]), 
         .Z(n14791)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6249_3_lut.init = 16'hcaca;
    LUT4 i5178_3_lut (.A(\array[62] [4]), .B(\array[63] [4]), .C(r_addr[0]), 
         .Z(n13720)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5178_3_lut.init = 16'hcaca;
    LUT4 i5177_3_lut (.A(\array[60] [4]), .B(\array[61] [4]), .C(r_addr[0]), 
         .Z(n13719)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5177_3_lut.init = 16'hcaca;
    LUT4 i5176_3_lut (.A(\array[58] [4]), .B(\array[59] [4]), .C(r_addr[0]), 
         .Z(n13718)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5176_3_lut.init = 16'hcaca;
    LUT4 i5175_3_lut (.A(\array[56] [4]), .B(\array[57] [4]), .C(r_addr[0]), 
         .Z(n13717)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5175_3_lut.init = 16'hcaca;
    LUT4 i5174_3_lut (.A(\array[54] [4]), .B(\array[55] [4]), .C(r_addr[0]), 
         .Z(n13716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5174_3_lut.init = 16'hcaca;
    LUT4 i5173_3_lut (.A(\array[52] [4]), .B(\array[53] [4]), .C(r_addr[0]), 
         .Z(n13715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5173_3_lut.init = 16'hcaca;
    LUT4 i5172_3_lut (.A(\array[50] [4]), .B(\array[51] [4]), .C(r_addr[0]), 
         .Z(n13714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5172_3_lut.init = 16'hcaca;
    LUT4 i5171_3_lut (.A(\array[48] [4]), .B(\array[49] [4]), .C(r_addr[0]), 
         .Z(n13713)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5171_3_lut.init = 16'hcaca;
    LUT4 i5170_3_lut (.A(\array[46] [4]), .B(\array[47] [4]), .C(r_addr[0]), 
         .Z(n13712)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5170_3_lut.init = 16'hcaca;
    LUT4 i5169_3_lut (.A(\array[44] [4]), .B(\array[45] [4]), .C(r_addr[0]), 
         .Z(n13711)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5169_3_lut.init = 16'hcaca;
    LUT4 i5168_3_lut (.A(\array[42] [4]), .B(\array[43] [4]), .C(r_addr[0]), 
         .Z(n13710)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5168_3_lut.init = 16'hcaca;
    LUT4 i5167_3_lut (.A(\array[40] [4]), .B(\array[41] [4]), .C(r_addr[0]), 
         .Z(n13709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5167_3_lut.init = 16'hcaca;
    LUT4 i5166_3_lut (.A(\array[38] [4]), .B(\array[39] [4]), .C(r_addr[0]), 
         .Z(n13708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5166_3_lut.init = 16'hcaca;
    LUT4 i4786_3_lut (.A(\array[178] [2]), .B(\array[179] [2]), .C(r_addr[0]), 
         .Z(n13328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4786_3_lut.init = 16'hcaca;
    LUT4 i4785_3_lut (.A(\array[176] [2]), .B(\array[177] [2]), .C(r_addr[0]), 
         .Z(n13327)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4785_3_lut.init = 16'hcaca;
    LUT4 i4784_3_lut (.A(\array[174] [2]), .B(\array[175] [2]), .C(r_addr[0]), 
         .Z(n13326)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4784_3_lut.init = 16'hcaca;
    LUT4 i4783_3_lut (.A(\array[172] [2]), .B(\array[173] [2]), .C(r_addr[0]), 
         .Z(n13325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4783_3_lut.init = 16'hcaca;
    LUT4 mux_4_i2_3_lut_4_lut (.A(n15023), .B(n15022), .C(\array[255] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_4097[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_4_i2_3_lut_4_lut.init = 16'hf870;
    LUT4 i4782_3_lut (.A(\array[170] [2]), .B(\array[171] [2]), .C(r_addr[0]), 
         .Z(n13324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4782_3_lut.init = 16'hcaca;
    LUT4 i4781_3_lut (.A(\array[168] [2]), .B(\array[169] [2]), .C(r_addr[0]), 
         .Z(n13323)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4781_3_lut.init = 16'hcaca;
    LUT4 i4780_3_lut (.A(\array[166] [2]), .B(\array[167] [2]), .C(r_addr[0]), 
         .Z(n13322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4780_3_lut.init = 16'hcaca;
    LUT4 i4779_3_lut (.A(\array[164] [2]), .B(\array[165] [2]), .C(r_addr[0]), 
         .Z(n13321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4779_3_lut.init = 16'hcaca;
    LUT4 i6001_3_lut (.A(\array[118] [7]), .B(\array[119] [7]), .C(r_addr[0]), 
         .Z(n14543)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6001_3_lut.init = 16'hcaca;
    LUT4 mux_4_i3_3_lut_4_lut (.A(n15023), .B(n15022), .C(\array[255] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_4097[2])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_4_i3_3_lut_4_lut.init = 16'hf870;
    LUT4 i6000_3_lut (.A(\array[116] [7]), .B(\array[117] [7]), .C(r_addr[0]), 
         .Z(n14542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6000_3_lut.init = 16'hcaca;
    LUT4 i4778_3_lut (.A(\array[162] [2]), .B(\array[163] [2]), .C(r_addr[0]), 
         .Z(n13320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4778_3_lut.init = 16'hcaca;
    LUT4 i4777_3_lut (.A(\array[160] [2]), .B(\array[161] [2]), .C(r_addr[0]), 
         .Z(n13319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4777_3_lut.init = 16'hcaca;
    LUT4 i5999_3_lut (.A(\array[114] [7]), .B(\array[115] [7]), .C(r_addr[0]), 
         .Z(n14541)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5999_3_lut.init = 16'hcaca;
    LUT4 mux_4_i4_3_lut_4_lut (.A(n15023), .B(n15022), .C(\array[255] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_4097[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_4_i4_3_lut_4_lut.init = 16'hf870;
    LUT4 i5998_3_lut (.A(\array[112] [7]), .B(\array[113] [7]), .C(r_addr[0]), 
         .Z(n14540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5998_3_lut.init = 16'hcaca;
    LUT4 i5997_3_lut (.A(\array[110] [7]), .B(\array[111] [7]), .C(r_addr[0]), 
         .Z(n14539)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5997_3_lut.init = 16'hcaca;
    LUT4 i5996_3_lut (.A(\array[108] [7]), .B(\array[109] [7]), .C(r_addr[0]), 
         .Z(n14538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5996_3_lut.init = 16'hcaca;
    LUT4 i5995_3_lut (.A(\array[106] [7]), .B(\array[107] [7]), .C(r_addr[0]), 
         .Z(n14537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5995_3_lut.init = 16'hcaca;
    LUT4 i5994_3_lut (.A(\array[104] [7]), .B(\array[105] [7]), .C(r_addr[0]), 
         .Z(n14536)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5994_3_lut.init = 16'hcaca;
    LUT4 mux_4_i5_3_lut_4_lut (.A(n15023), .B(n15022), .C(\array[255] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_4097[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_4_i5_3_lut_4_lut.init = 16'hf870;
    LUT4 i5993_3_lut (.A(\array[102] [7]), .B(\array[103] [7]), .C(r_addr[0]), 
         .Z(n14535)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5993_3_lut.init = 16'hcaca;
    LUT4 i5992_3_lut (.A(\array[100] [7]), .B(\array[101] [7]), .C(r_addr[0]), 
         .Z(n14534)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5992_3_lut.init = 16'hcaca;
    LUT4 i5588_3_lut (.A(\array[222] [5]), .B(\array[223] [5]), .C(r_addr[0]), 
         .Z(n14130)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5588_3_lut.init = 16'hcaca;
    LUT4 i5587_3_lut (.A(\array[220] [5]), .B(\array[221] [5]), .C(r_addr[0]), 
         .Z(n14129)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5587_3_lut.init = 16'hcaca;
    LUT4 i5991_3_lut (.A(\array[98] [7]), .B(\array[99] [7]), .C(r_addr[0]), 
         .Z(n14533)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5991_3_lut.init = 16'hcaca;
    LUT4 mux_4_i6_3_lut_4_lut (.A(n15023), .B(n15022), .C(\array[255] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_4097[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_4_i6_3_lut_4_lut.init = 16'hf870;
    LUT4 i5990_3_lut (.A(\array[96] [7]), .B(\array[97] [7]), .C(r_addr[0]), 
         .Z(n14532)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5990_3_lut.init = 16'hcaca;
    LUT4 i5586_3_lut (.A(\array[218] [5]), .B(\array[219] [5]), .C(r_addr[0]), 
         .Z(n14128)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5586_3_lut.init = 16'hcaca;
    LUT4 i5585_3_lut (.A(\array[216] [5]), .B(\array[217] [5]), .C(r_addr[0]), 
         .Z(n14127)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5585_3_lut.init = 16'hcaca;
    LUT4 i4761_3_lut (.A(\array[158] [2]), .B(\array[159] [2]), .C(r_addr[0]), 
         .Z(n13303)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4761_3_lut.init = 16'hcaca;
    LUT4 i4760_3_lut (.A(\array[156] [2]), .B(\array[157] [2]), .C(r_addr[0]), 
         .Z(n13302)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4760_3_lut.init = 16'hcaca;
    LUT4 mux_4_i7_3_lut_4_lut (.A(n15023), .B(n15022), .C(\array[255] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_4097[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_4_i7_3_lut_4_lut.init = 16'hf870;
    LUT4 i5584_3_lut (.A(\array[214] [5]), .B(\array[215] [5]), .C(r_addr[0]), 
         .Z(n14126)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5584_3_lut.init = 16'hcaca;
    LUT4 i5583_3_lut (.A(\array[212] [5]), .B(\array[213] [5]), .C(r_addr[0]), 
         .Z(n14125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5583_3_lut.init = 16'hcaca;
    LUT4 i4759_3_lut (.A(\array[154] [2]), .B(\array[155] [2]), .C(r_addr[0]), 
         .Z(n13301)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4759_3_lut.init = 16'hcaca;
    LUT4 i4758_3_lut (.A(\array[152] [2]), .B(\array[153] [2]), .C(r_addr[0]), 
         .Z(n13300)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4758_3_lut.init = 16'hcaca;
    LUT4 i4757_3_lut (.A(\array[150] [2]), .B(\array[151] [2]), .C(r_addr[0]), 
         .Z(n13299)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4757_3_lut.init = 16'hcaca;
    LUT4 mux_4_i8_3_lut_4_lut (.A(n15023), .B(n15022), .C(\array[255] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_4097[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_4_i8_3_lut_4_lut.init = 16'hf870;
    LUT4 i4756_3_lut (.A(\array[148] [2]), .B(\array[149] [2]), .C(r_addr[0]), 
         .Z(n13298)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4756_3_lut.init = 16'hcaca;
    LUT4 i5582_3_lut (.A(\array[210] [5]), .B(\array[211] [5]), .C(r_addr[0]), 
         .Z(n14124)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5582_3_lut.init = 16'hcaca;
    LUT4 i5581_3_lut (.A(\array[208] [5]), .B(\array[209] [5]), .C(r_addr[0]), 
         .Z(n14123)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5581_3_lut.init = 16'hcaca;
    LUT4 i4755_3_lut (.A(\array[146] [2]), .B(\array[147] [2]), .C(r_addr[0]), 
         .Z(n13297)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4755_3_lut.init = 16'hcaca;
    LUT4 i4754_3_lut (.A(\array[144] [2]), .B(\array[145] [2]), .C(r_addr[0]), 
         .Z(n13296)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4754_3_lut.init = 16'hcaca;
    LUT4 i4753_3_lut (.A(\array[142] [2]), .B(\array[143] [2]), .C(r_addr[0]), 
         .Z(n13295)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4753_3_lut.init = 16'hcaca;
    LUT4 i4752_3_lut (.A(\array[140] [2]), .B(\array[141] [2]), .C(r_addr[0]), 
         .Z(n13294)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4752_3_lut.init = 16'hcaca;
    LUT4 i5580_3_lut (.A(\array[206] [5]), .B(\array[207] [5]), .C(r_addr[0]), 
         .Z(n14122)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5580_3_lut.init = 16'hcaca;
    LUT4 mux_253_i2_3_lut_4_lut (.A(n15013), .B(n14992), .C(\array[6] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2105[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_253_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5579_3_lut (.A(\array[204] [5]), .B(\array[205] [5]), .C(r_addr[0]), 
         .Z(n14121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5579_3_lut.init = 16'hcaca;
    LUT4 i4751_3_lut (.A(\array[138] [2]), .B(\array[139] [2]), .C(r_addr[0]), 
         .Z(n13293)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4751_3_lut.init = 16'hcaca;
    LUT4 i4750_3_lut (.A(\array[136] [2]), .B(\array[137] [2]), .C(r_addr[0]), 
         .Z(n13292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4750_3_lut.init = 16'hcaca;
    LUT4 i4749_3_lut (.A(\array[134] [2]), .B(\array[135] [2]), .C(r_addr[0]), 
         .Z(n13291)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4749_3_lut.init = 16'hcaca;
    LUT4 i4748_3_lut (.A(\array[132] [2]), .B(\array[133] [2]), .C(r_addr[0]), 
         .Z(n13290)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4748_3_lut.init = 16'hcaca;
    LUT4 i5578_3_lut (.A(\array[202] [5]), .B(\array[203] [5]), .C(r_addr[0]), 
         .Z(n14120)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5578_3_lut.init = 16'hcaca;
    LUT4 i5577_3_lut (.A(\array[200] [5]), .B(\array[201] [5]), .C(r_addr[0]), 
         .Z(n14119)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5577_3_lut.init = 16'hcaca;
    LUT4 i4747_3_lut (.A(\array[130] [2]), .B(\array[131] [2]), .C(r_addr[0]), 
         .Z(n13289)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4747_3_lut.init = 16'hcaca;
    LUT4 mux_253_i3_3_lut_4_lut (.A(n15013), .B(n14992), .C(\array[6] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2105[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_253_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4746_3_lut (.A(\array[128] [2]), .B(\array[129] [2]), .C(r_addr[0]), 
         .Z(n13288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4746_3_lut.init = 16'hcaca;
    LUT4 i5576_3_lut (.A(\array[198] [5]), .B(\array[199] [5]), .C(r_addr[0]), 
         .Z(n14118)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5576_3_lut.init = 16'hcaca;
    LUT4 i5575_3_lut (.A(\array[196] [5]), .B(\array[197] [5]), .C(r_addr[0]), 
         .Z(n14117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5575_3_lut.init = 16'hcaca;
    LUT4 i6380_3_lut (.A(\array[246] [0]), .B(\array[247] [0]), .C(r_addr[0]), 
         .Z(n14922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6380_3_lut.init = 16'hcaca;
    LUT4 i6379_3_lut (.A(\array[244] [0]), .B(\array[245] [0]), .C(r_addr[0]), 
         .Z(n14921)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6379_3_lut.init = 16'hcaca;
    LUT4 i5574_3_lut (.A(\array[194] [5]), .B(\array[195] [5]), .C(r_addr[0]), 
         .Z(n14116)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5574_3_lut.init = 16'hcaca;
    LUT4 i5573_3_lut (.A(\array[192] [5]), .B(\array[193] [5]), .C(r_addr[0]), 
         .Z(n14115)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5573_3_lut.init = 16'hcaca;
    LUT4 i4730_3_lut (.A(\array[126] [2]), .B(\array[127] [2]), .C(r_addr[0]), 
         .Z(n13272)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4730_3_lut.init = 16'hcaca;
    VHI i4126 (.Z(VCC_net));
    LUT4 i4729_3_lut (.A(\array[124] [2]), .B(\array[125] [2]), .C(r_addr[0]), 
         .Z(n13271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4729_3_lut.init = 16'hcaca;
    LUT4 i4728_3_lut (.A(\array[122] [2]), .B(\array[123] [2]), .C(r_addr[0]), 
         .Z(n13270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4728_3_lut.init = 16'hcaca;
    LUT4 i4727_3_lut (.A(\array[120] [2]), .B(\array[121] [2]), .C(r_addr[0]), 
         .Z(n13269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4727_3_lut.init = 16'hcaca;
    LUT4 i4726_3_lut (.A(\array[118] [2]), .B(\array[119] [2]), .C(r_addr[0]), 
         .Z(n13268)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4726_3_lut.init = 16'hcaca;
    LUT4 i4725_3_lut (.A(\array[116] [2]), .B(\array[117] [2]), .C(r_addr[0]), 
         .Z(n13267)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4725_3_lut.init = 16'hcaca;
    TSALL TSALL_INST (.TSALL(GND_net));
    LUT4 i6198_3_lut (.A(\array[62] [0]), .B(\array[63] [0]), .C(r_addr[0]), 
         .Z(n14740)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6198_3_lut.init = 16'hcaca;
    LUT4 i6197_3_lut (.A(\array[60] [0]), .B(\array[61] [0]), .C(r_addr[0]), 
         .Z(n14739)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6197_3_lut.init = 16'hcaca;
    LUT4 i4724_3_lut (.A(\array[114] [2]), .B(\array[115] [2]), .C(r_addr[0]), 
         .Z(n13266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4724_3_lut.init = 16'hcaca;
    LUT4 i4723_3_lut (.A(\array[112] [2]), .B(\array[113] [2]), .C(r_addr[0]), 
         .Z(n13265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4723_3_lut.init = 16'hcaca;
    LUT4 i4722_3_lut (.A(\array[110] [2]), .B(\array[111] [2]), .C(r_addr[0]), 
         .Z(n13264)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4722_3_lut.init = 16'hcaca;
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i4721_3_lut (.A(\array[108] [2]), .B(\array[109] [2]), .C(r_addr[0]), 
         .Z(n13263)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4721_3_lut.init = 16'hcaca;
    LUT4 i4720_3_lut (.A(\array[106] [2]), .B(\array[107] [2]), .C(r_addr[0]), 
         .Z(n13262)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4720_3_lut.init = 16'hcaca;
    LUT4 i4719_3_lut (.A(\array[104] [2]), .B(\array[105] [2]), .C(r_addr[0]), 
         .Z(n13261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4719_3_lut.init = 16'hcaca;
    LUT4 i4718_3_lut (.A(\array[102] [2]), .B(\array[103] [2]), .C(r_addr[0]), 
         .Z(n13260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4718_3_lut.init = 16'hcaca;
    LUT4 i4717_3_lut (.A(\array[100] [2]), .B(\array[101] [2]), .C(r_addr[0]), 
         .Z(n13259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4717_3_lut.init = 16'hcaca;
    FD1P3AX r_addr_i0_i0_rep_92 (.D(addr_c_0), .SP(clk_c_enable_2057), .CK(clk_c), 
            .Q(maxfan_replicated_net_23)) /* synthesis maxfan_replicated_inst=1 */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam r_addr_i0_i0_rep_92.GSR = "ENABLED";
    LUT4 i4716_3_lut (.A(\array[98] [2]), .B(\array[99] [2]), .C(r_addr[0]), 
         .Z(n13258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4716_3_lut.init = 16'hcaca;
    LUT4 i4715_3_lut (.A(\array[96] [2]), .B(\array[97] [2]), .C(r_addr[0]), 
         .Z(n13257)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4715_3_lut.init = 16'hcaca;
    LUT4 i6196_3_lut (.A(\array[58] [0]), .B(\array[59] [0]), .C(r_addr[0]), 
         .Z(n14738)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6196_3_lut.init = 16'hcaca;
    LUT4 i6195_3_lut (.A(\array[56] [0]), .B(\array[57] [0]), .C(r_addr[0]), 
         .Z(n14737)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6195_3_lut.init = 16'hcaca;
    LUT4 i6194_3_lut (.A(\array[54] [0]), .B(\array[55] [0]), .C(r_addr[0]), 
         .Z(n14736)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6194_3_lut.init = 16'hcaca;
    LUT4 i6193_3_lut (.A(\array[52] [0]), .B(\array[53] [0]), .C(r_addr[0]), 
         .Z(n14735)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6193_3_lut.init = 16'hcaca;
    LUT4 i5557_3_lut (.A(\array[190] [5]), .B(\array[191] [5]), .C(r_addr[0]), 
         .Z(n14099)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5557_3_lut.init = 16'hcaca;
    LUT4 i5556_3_lut (.A(\array[188] [5]), .B(\array[189] [5]), .C(r_addr[0]), 
         .Z(n14098)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5556_3_lut.init = 16'hcaca;
    LUT4 i6192_3_lut (.A(\array[50] [0]), .B(\array[51] [0]), .C(r_addr[0]), 
         .Z(n14734)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6192_3_lut.init = 16'hcaca;
    LUT4 i6191_3_lut (.A(\array[48] [0]), .B(\array[49] [0]), .C(r_addr[0]), 
         .Z(n14733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6191_3_lut.init = 16'hcaca;
    LUT4 i5555_3_lut (.A(\array[186] [5]), .B(\array[187] [5]), .C(r_addr[0]), 
         .Z(n14097)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5555_3_lut.init = 16'hcaca;
    LUT4 i5554_3_lut (.A(\array[184] [5]), .B(\array[185] [5]), .C(r_addr[0]), 
         .Z(n14096)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5554_3_lut.init = 16'hcaca;
    LUT4 i4699_3_lut (.A(\array[94] [2]), .B(\array[95] [2]), .C(r_addr[0]), 
         .Z(n13241)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4699_3_lut.init = 16'hcaca;
    LUT4 i4698_3_lut (.A(\array[92] [2]), .B(\array[93] [2]), .C(r_addr[0]), 
         .Z(n13240)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4698_3_lut.init = 16'hcaca;
    LUT4 i5553_3_lut (.A(\array[182] [5]), .B(\array[183] [5]), .C(r_addr[0]), 
         .Z(n14095)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5553_3_lut.init = 16'hcaca;
    LUT4 i5552_3_lut (.A(\array[180] [5]), .B(\array[181] [5]), .C(r_addr[0]), 
         .Z(n14094)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5552_3_lut.init = 16'hcaca;
    LUT4 i4697_3_lut (.A(\array[90] [2]), .B(\array[91] [2]), .C(r_addr[0]), 
         .Z(n13239)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4697_3_lut.init = 16'hcaca;
    LUT4 i4696_3_lut (.A(\array[88] [2]), .B(\array[89] [2]), .C(r_addr[0]), 
         .Z(n13238)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4696_3_lut.init = 16'hcaca;
    LUT4 i4695_3_lut (.A(\array[86] [2]), .B(\array[87] [2]), .C(r_addr[0]), 
         .Z(n13237)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4695_3_lut.init = 16'hcaca;
    LUT4 i4694_3_lut (.A(\array[84] [2]), .B(\array[85] [2]), .C(r_addr[0]), 
         .Z(n13236)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4694_3_lut.init = 16'hcaca;
    LUT4 i5551_3_lut (.A(\array[178] [5]), .B(\array[179] [5]), .C(r_addr[0]), 
         .Z(n14093)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5551_3_lut.init = 16'hcaca;
    LUT4 i5550_3_lut (.A(\array[176] [5]), .B(\array[177] [5]), .C(r_addr[0]), 
         .Z(n14092)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5550_3_lut.init = 16'hcaca;
    LUT4 i4693_3_lut (.A(\array[82] [2]), .B(\array[83] [2]), .C(r_addr[0]), 
         .Z(n13235)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4693_3_lut.init = 16'hcaca;
    LUT4 i4692_3_lut (.A(\array[80] [2]), .B(\array[81] [2]), .C(r_addr[0]), 
         .Z(n13234)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4692_3_lut.init = 16'hcaca;
    LUT4 i4691_3_lut (.A(\array[78] [2]), .B(\array[79] [2]), .C(r_addr[0]), 
         .Z(n13233)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4691_3_lut.init = 16'hcaca;
    LUT4 i4690_3_lut (.A(\array[76] [2]), .B(\array[77] [2]), .C(r_addr[0]), 
         .Z(n13232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4690_3_lut.init = 16'hcaca;
    LUT4 i5549_3_lut (.A(\array[174] [5]), .B(\array[175] [5]), .C(r_addr[0]), 
         .Z(n14091)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5549_3_lut.init = 16'hcaca;
    LUT4 i5548_3_lut (.A(\array[172] [5]), .B(\array[173] [5]), .C(r_addr[0]), 
         .Z(n14090)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5548_3_lut.init = 16'hcaca;
    LUT4 i6190_3_lut (.A(\array[46] [0]), .B(\array[47] [0]), .C(r_addr[0]), 
         .Z(n14732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6190_3_lut.init = 16'hcaca;
    LUT4 i6189_3_lut (.A(\array[44] [0]), .B(\array[45] [0]), .C(r_addr[0]), 
         .Z(n14731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6189_3_lut.init = 16'hcaca;
    LUT4 i4689_3_lut (.A(\array[74] [2]), .B(\array[75] [2]), .C(r_addr[0]), 
         .Z(n13231)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4689_3_lut.init = 16'hcaca;
    LUT4 i4688_3_lut (.A(\array[72] [2]), .B(\array[73] [2]), .C(r_addr[0]), 
         .Z(n13230)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4688_3_lut.init = 16'hcaca;
    LUT4 i4687_3_lut (.A(\array[70] [2]), .B(\array[71] [2]), .C(r_addr[0]), 
         .Z(n13229)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4687_3_lut.init = 16'hcaca;
    LUT4 i4686_3_lut (.A(\array[68] [2]), .B(\array[69] [2]), .C(r_addr[0]), 
         .Z(n13228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4686_3_lut.init = 16'hcaca;
    LUT4 i5547_3_lut (.A(\array[170] [5]), .B(\array[171] [5]), .C(r_addr[0]), 
         .Z(n14089)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5547_3_lut.init = 16'hcaca;
    LUT4 i5546_3_lut (.A(\array[168] [5]), .B(\array[169] [5]), .C(r_addr[0]), 
         .Z(n14088)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5546_3_lut.init = 16'hcaca;
    LUT4 i4685_3_lut (.A(\array[66] [2]), .B(\array[67] [2]), .C(r_addr[0]), 
         .Z(n13227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4685_3_lut.init = 16'hcaca;
    LUT4 i4684_3_lut (.A(\array[64] [2]), .B(\array[65] [2]), .C(r_addr[0]), 
         .Z(n13226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4684_3_lut.init = 16'hcaca;
    LUT4 i5545_3_lut (.A(\array[166] [5]), .B(\array[167] [5]), .C(r_addr[0]), 
         .Z(n14087)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5545_3_lut.init = 16'hcaca;
    LUT4 i5544_3_lut (.A(\array[164] [5]), .B(\array[165] [5]), .C(r_addr[0]), 
         .Z(n14086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5544_3_lut.init = 16'hcaca;
    LUT4 i5543_3_lut (.A(\array[162] [5]), .B(\array[163] [5]), .C(r_addr[0]), 
         .Z(n14085)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5543_3_lut.init = 16'hcaca;
    LUT4 i5542_3_lut (.A(\array[160] [5]), .B(\array[161] [5]), .C(r_addr[0]), 
         .Z(n14084)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5542_3_lut.init = 16'hcaca;
    LUT4 i6188_3_lut (.A(\array[42] [0]), .B(\array[43] [0]), .C(r_addr[0]), 
         .Z(n14730)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6188_3_lut.init = 16'hcaca;
    LUT4 i6187_3_lut (.A(\array[40] [0]), .B(\array[41] [0]), .C(r_addr[0]), 
         .Z(n14729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6187_3_lut.init = 16'hcaca;
    LUT4 i6378_3_lut (.A(\array[242] [0]), .B(\array[243] [0]), .C(r_addr[0]), 
         .Z(n14920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6378_3_lut.init = 16'hcaca;
    LUT4 i6377_3_lut (.A(\array[240] [0]), .B(\array[241] [0]), .C(r_addr[0]), 
         .Z(n14919)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6377_3_lut.init = 16'hcaca;
    LUT4 i6186_3_lut (.A(\array[38] [0]), .B(\array[39] [0]), .C(r_addr[0]), 
         .Z(n14728)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6186_3_lut.init = 16'hcaca;
    LUT4 i6185_3_lut (.A(\array[36] [0]), .B(\array[37] [0]), .C(r_addr[0]), 
         .Z(n14727)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6185_3_lut.init = 16'hcaca;
    LUT4 i5974_3_lut (.A(\array[94] [7]), .B(\array[95] [7]), .C(r_addr[0]), 
         .Z(n14516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5974_3_lut.init = 16'hcaca;
    LUT4 i5973_3_lut (.A(\array[92] [7]), .B(\array[93] [7]), .C(r_addr[0]), 
         .Z(n14515)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5973_3_lut.init = 16'hcaca;
    LUT4 i6184_3_lut (.A(\array[34] [0]), .B(\array[35] [0]), .C(r_addr[0]), 
         .Z(n14726)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6184_3_lut.init = 16'hcaca;
    LUT4 i6183_3_lut (.A(\array[32] [0]), .B(\array[33] [0]), .C(r_addr[0]), 
         .Z(n14725)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6183_3_lut.init = 16'hcaca;
    LUT4 i4668_3_lut (.A(\array[62] [2]), .B(\array[63] [2]), .C(r_addr[0]), 
         .Z(n13210)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4668_3_lut.init = 16'hcaca;
    LUT4 i4667_3_lut (.A(\array[60] [2]), .B(\array[61] [2]), .C(r_addr[0]), 
         .Z(n13209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4667_3_lut.init = 16'hcaca;
    LUT4 i4666_3_lut (.A(\array[58] [2]), .B(\array[59] [2]), .C(r_addr[0]), 
         .Z(n13208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4666_3_lut.init = 16'hcaca;
    LUT4 i4665_3_lut (.A(\array[56] [2]), .B(\array[57] [2]), .C(r_addr[0]), 
         .Z(n13207)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4665_3_lut.init = 16'hcaca;
    LUT4 i5972_3_lut (.A(\array[90] [7]), .B(\array[91] [7]), .C(r_addr[0]), 
         .Z(n14514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5972_3_lut.init = 16'hcaca;
    LUT4 i5971_3_lut (.A(\array[88] [7]), .B(\array[89] [7]), .C(r_addr[0]), 
         .Z(n14513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5971_3_lut.init = 16'hcaca;
    LUT4 i4664_3_lut (.A(\array[54] [2]), .B(\array[55] [2]), .C(r_addr[0]), 
         .Z(n13206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4664_3_lut.init = 16'hcaca;
    LUT4 i4663_3_lut (.A(\array[52] [2]), .B(\array[53] [2]), .C(r_addr[0]), 
         .Z(n13205)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4663_3_lut.init = 16'hcaca;
    LUT4 i4662_3_lut (.A(\array[50] [2]), .B(\array[51] [2]), .C(r_addr[0]), 
         .Z(n13204)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4662_3_lut.init = 16'hcaca;
    LUT4 i4661_3_lut (.A(\array[48] [2]), .B(\array[49] [2]), .C(r_addr[0]), 
         .Z(n13203)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4661_3_lut.init = 16'hcaca;
    LUT4 i4660_3_lut (.A(\array[46] [2]), .B(\array[47] [2]), .C(r_addr[0]), 
         .Z(n13202)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4660_3_lut.init = 16'hcaca;
    LUT4 i4659_3_lut (.A(\array[44] [2]), .B(\array[45] [2]), .C(r_addr[0]), 
         .Z(n13201)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4659_3_lut.init = 16'hcaca;
    LUT4 i4658_3_lut (.A(\array[42] [2]), .B(\array[43] [2]), .C(r_addr[0]), 
         .Z(n13200)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4658_3_lut.init = 16'hcaca;
    LUT4 i4657_3_lut (.A(\array[40] [2]), .B(\array[41] [2]), .C(r_addr[0]), 
         .Z(n13199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4657_3_lut.init = 16'hcaca;
    LUT4 i5970_3_lut (.A(\array[86] [7]), .B(\array[87] [7]), .C(r_addr[0]), 
         .Z(n14512)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5970_3_lut.init = 16'hcaca;
    LUT4 i5969_3_lut (.A(\array[84] [7]), .B(\array[85] [7]), .C(r_addr[0]), 
         .Z(n14511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5969_3_lut.init = 16'hcaca;
    LUT4 i4656_3_lut (.A(\array[38] [2]), .B(\array[39] [2]), .C(r_addr[0]), 
         .Z(n13198)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4656_3_lut.init = 16'hcaca;
    LUT4 i4655_3_lut (.A(\array[36] [2]), .B(\array[37] [2]), .C(r_addr[0]), 
         .Z(n13197)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4655_3_lut.init = 16'hcaca;
    LUT4 i4654_3_lut (.A(\array[34] [2]), .B(\array[35] [2]), .C(r_addr[0]), 
         .Z(n13196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4654_3_lut.init = 16'hcaca;
    LUT4 i4653_3_lut (.A(\array[32] [2]), .B(\array[33] [2]), .C(r_addr[0]), 
         .Z(n13195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4653_3_lut.init = 16'hcaca;
    LUT4 i5968_3_lut (.A(\array[82] [7]), .B(\array[83] [7]), .C(r_addr[0]), 
         .Z(n14510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5968_3_lut.init = 16'hcaca;
    LUT4 i5967_3_lut (.A(\array[80] [7]), .B(\array[81] [7]), .C(r_addr[0]), 
         .Z(n14509)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5967_3_lut.init = 16'hcaca;
    LUT4 i5966_3_lut (.A(\array[78] [7]), .B(\array[79] [7]), .C(r_addr[0]), 
         .Z(n14508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5966_3_lut.init = 16'hcaca;
    LUT4 i5965_3_lut (.A(\array[76] [7]), .B(\array[77] [7]), .C(r_addr[0]), 
         .Z(n14507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5965_3_lut.init = 16'hcaca;
    LUT4 i6353_3_lut (.A(\array[222] [0]), .B(\array[223] [0]), .C(r_addr[0]), 
         .Z(n14895)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6353_3_lut.init = 16'hcaca;
    LUT4 i6352_3_lut (.A(\array[220] [0]), .B(\array[221] [0]), .C(r_addr[0]), 
         .Z(n14894)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6352_3_lut.init = 16'hcaca;
    LUT4 i5964_3_lut (.A(\array[74] [7]), .B(\array[75] [7]), .C(r_addr[0]), 
         .Z(n14506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5964_3_lut.init = 16'hcaca;
    LUT4 i5963_3_lut (.A(\array[72] [7]), .B(\array[73] [7]), .C(r_addr[0]), 
         .Z(n14505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5963_3_lut.init = 16'hcaca;
    LUT4 i5962_3_lut (.A(\array[70] [7]), .B(\array[71] [7]), .C(r_addr[0]), 
         .Z(n14504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5962_3_lut.init = 16'hcaca;
    LUT4 i5961_3_lut (.A(\array[68] [7]), .B(\array[69] [7]), .C(r_addr[0]), 
         .Z(n14503)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5961_3_lut.init = 16'hcaca;
    LUT4 i5526_3_lut (.A(\array[158] [5]), .B(\array[159] [5]), .C(r_addr[0]), 
         .Z(n14068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5526_3_lut.init = 16'hcaca;
    LUT4 i5525_3_lut (.A(\array[156] [5]), .B(\array[157] [5]), .C(r_addr[0]), 
         .Z(n14067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5525_3_lut.init = 16'hcaca;
    LUT4 i5960_3_lut (.A(\array[66] [7]), .B(\array[67] [7]), .C(r_addr[0]), 
         .Z(n14502)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5960_3_lut.init = 16'hcaca;
    LUT4 i5959_3_lut (.A(\array[64] [7]), .B(\array[65] [7]), .C(r_addr[0]), 
         .Z(n14501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5959_3_lut.init = 16'hcaca;
    LUT4 i5524_3_lut (.A(\array[154] [5]), .B(\array[155] [5]), .C(r_addr[0]), 
         .Z(n14066)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5524_3_lut.init = 16'hcaca;
    LUT4 i5523_3_lut (.A(\array[152] [5]), .B(\array[153] [5]), .C(r_addr[0]), 
         .Z(n14065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5523_3_lut.init = 16'hcaca;
    LUT4 i5522_3_lut (.A(\array[150] [5]), .B(\array[151] [5]), .C(r_addr[0]), 
         .Z(n14064)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5522_3_lut.init = 16'hcaca;
    LUT4 i5521_3_lut (.A(\array[148] [5]), .B(\array[149] [5]), .C(r_addr[0]), 
         .Z(n14063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5521_3_lut.init = 16'hcaca;
    LUT4 i4637_3_lut (.A(\array[30] [2]), .B(\array[31] [2]), .C(r_addr[0]), 
         .Z(n13179)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4637_3_lut.init = 16'hcaca;
    LUT4 i4636_3_lut (.A(\array[28] [2]), .B(\array[29] [2]), .C(r_addr[0]), 
         .Z(n13178)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4636_3_lut.init = 16'hcaca;
    LUT4 i4635_3_lut (.A(\array[26] [2]), .B(\array[27] [2]), .C(r_addr[0]), 
         .Z(n13177)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4635_3_lut.init = 16'hcaca;
    LUT4 i4634_3_lut (.A(\array[24] [2]), .B(\array[25] [2]), .C(r_addr[0]), 
         .Z(n13176)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4634_3_lut.init = 16'hcaca;
    LUT4 i5520_3_lut (.A(\array[146] [5]), .B(\array[147] [5]), .C(r_addr[0]), 
         .Z(n14062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5520_3_lut.init = 16'hcaca;
    LUT4 i5519_3_lut (.A(\array[144] [5]), .B(\array[145] [5]), .C(r_addr[0]), 
         .Z(n14061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5519_3_lut.init = 16'hcaca;
    LUT4 i4633_3_lut (.A(\array[22] [2]), .B(\array[23] [2]), .C(r_addr[0]), 
         .Z(n13175)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4633_3_lut.init = 16'hcaca;
    LUT4 i4632_3_lut (.A(\array[20] [2]), .B(\array[21] [2]), .C(r_addr[0]), 
         .Z(n13174)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4632_3_lut.init = 16'hcaca;
    LUT4 i4631_3_lut (.A(\array[18] [2]), .B(\array[19] [2]), .C(r_addr[0]), 
         .Z(n13173)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4631_3_lut.init = 16'hcaca;
    LUT4 i4630_3_lut (.A(\array[16] [2]), .B(\array[17] [2]), .C(r_addr[0]), 
         .Z(n13172)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4630_3_lut.init = 16'hcaca;
    LUT4 i5518_3_lut (.A(\array[142] [5]), .B(\array[143] [5]), .C(r_addr[0]), 
         .Z(n14060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5518_3_lut.init = 16'hcaca;
    LUT4 i5517_3_lut (.A(\array[140] [5]), .B(\array[141] [5]), .C(r_addr[0]), 
         .Z(n14059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5517_3_lut.init = 16'hcaca;
    LUT4 i4629_3_lut (.A(\array[14] [2]), .B(\array[15] [2]), .C(r_addr[0]), 
         .Z(n13171)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4629_3_lut.init = 16'hcaca;
    LUT4 i4628_3_lut (.A(\array[12] [2]), .B(\array[13] [2]), .C(r_addr[0]), 
         .Z(n13170)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4628_3_lut.init = 16'hcaca;
    LUT4 i4627_3_lut (.A(\array[10] [2]), .B(\array[11] [2]), .C(r_addr[0]), 
         .Z(n13169)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4627_3_lut.init = 16'hcaca;
    LUT4 i4626_3_lut (.A(\array[8] [2]), .B(\array[9] [2]), .C(r_addr[0]), 
         .Z(n13168)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4626_3_lut.init = 16'hcaca;
    LUT4 i5516_3_lut (.A(\array[138] [5]), .B(\array[139] [5]), .C(r_addr[0]), 
         .Z(n14058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5516_3_lut.init = 16'hcaca;
    LUT4 i5515_3_lut (.A(\array[136] [5]), .B(\array[137] [5]), .C(r_addr[0]), 
         .Z(n14057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5515_3_lut.init = 16'hcaca;
    LUT4 i4625_3_lut (.A(\array[6] [2]), .B(\array[7] [2]), .C(r_addr[0]), 
         .Z(n13167)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4625_3_lut.init = 16'hcaca;
    LUT4 i4624_3_lut (.A(\array[4] [2]), .B(\array[5] [2]), .C(r_addr[0]), 
         .Z(n13166)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4624_3_lut.init = 16'hcaca;
    LUT4 i4623_3_lut (.A(\array[2] [2]), .B(\array[3] [2]), .C(r_addr[0]), 
         .Z(n13165)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4623_3_lut.init = 16'hcaca;
    LUT4 i4622_3_lut (.A(\array[0] [2]), .B(\array[1] [2]), .C(r_addr[0]), 
         .Z(n13164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4622_3_lut.init = 16'hcaca;
    LUT4 i5514_3_lut (.A(\array[134] [5]), .B(\array[135] [5]), .C(r_addr[0]), 
         .Z(n14056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5514_3_lut.init = 16'hcaca;
    LUT4 i5513_3_lut (.A(\array[132] [5]), .B(\array[133] [5]), .C(r_addr[0]), 
         .Z(n14055)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5513_3_lut.init = 16'hcaca;
    LUT4 i5512_3_lut (.A(\array[130] [5]), .B(\array[131] [5]), .C(r_addr[0]), 
         .Z(n14054)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5512_3_lut.init = 16'hcaca;
    LUT4 i5511_3_lut (.A(\array[128] [5]), .B(\array[129] [5]), .C(r_addr[0]), 
         .Z(n14053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5511_3_lut.init = 16'hcaca;
    LUT4 i6351_3_lut (.A(\array[218] [0]), .B(\array[219] [0]), .C(r_addr[0]), 
         .Z(n14893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6351_3_lut.init = 16'hcaca;
    LUT4 i6350_3_lut (.A(\array[216] [0]), .B(\array[217] [0]), .C(r_addr[0]), 
         .Z(n14892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6350_3_lut.init = 16'hcaca;
    LUT4 i6376_3_lut (.A(\array[238] [0]), .B(\array[239] [0]), .C(r_addr[0]), 
         .Z(n14918)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6376_3_lut.init = 16'hcaca;
    LUT4 i6375_3_lut (.A(\array[236] [0]), .B(\array[237] [0]), .C(r_addr[0]), 
         .Z(n14917)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6375_3_lut.init = 16'hcaca;
    LUT4 i4599_3_lut (.A(\array[254] [1]), .B(\array[255] [1]), .C(r_addr[0]), 
         .Z(n13141)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4599_3_lut.init = 16'hcaca;
    LUT4 i4598_3_lut (.A(\array[252] [1]), .B(\array[253] [1]), .C(r_addr[0]), 
         .Z(n13140)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4598_3_lut.init = 16'hcaca;
    LUT4 i4597_3_lut (.A(\array[250] [1]), .B(\array[251] [1]), .C(r_addr[0]), 
         .Z(n13139)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4597_3_lut.init = 16'hcaca;
    LUT4 i4596_3_lut (.A(\array[248] [1]), .B(\array[249] [1]), .C(r_addr[0]), 
         .Z(n13138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4596_3_lut.init = 16'hcaca;
    LUT4 i4595_3_lut (.A(\array[246] [1]), .B(\array[247] [1]), .C(r_addr[0]), 
         .Z(n13137)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4595_3_lut.init = 16'hcaca;
    LUT4 i4594_3_lut (.A(\array[244] [1]), .B(\array[245] [1]), .C(r_addr[0]), 
         .Z(n13136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4594_3_lut.init = 16'hcaca;
    LUT4 i4593_3_lut (.A(\array[242] [1]), .B(\array[243] [1]), .C(r_addr[0]), 
         .Z(n13135)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4593_3_lut.init = 16'hcaca;
    LUT4 i4592_3_lut (.A(\array[240] [1]), .B(\array[241] [1]), .C(r_addr[0]), 
         .Z(n13134)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4592_3_lut.init = 16'hcaca;
    LUT4 i4591_3_lut (.A(\array[238] [1]), .B(\array[239] [1]), .C(r_addr[0]), 
         .Z(n13133)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4591_3_lut.init = 16'hcaca;
    LUT4 i4590_3_lut (.A(\array[236] [1]), .B(\array[237] [1]), .C(r_addr[0]), 
         .Z(n13132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4590_3_lut.init = 16'hcaca;
    LUT4 i4589_3_lut (.A(\array[234] [1]), .B(\array[235] [1]), .C(r_addr[0]), 
         .Z(n13131)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4589_3_lut.init = 16'hcaca;
    LUT4 i4588_3_lut (.A(\array[232] [1]), .B(\array[233] [1]), .C(r_addr[0]), 
         .Z(n13130)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4588_3_lut.init = 16'hcaca;
    LUT4 i4587_3_lut (.A(\array[230] [1]), .B(\array[231] [1]), .C(r_addr[0]), 
         .Z(n13129)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4587_3_lut.init = 16'hcaca;
    LUT4 i4586_3_lut (.A(\array[228] [1]), .B(\array[229] [1]), .C(r_addr[0]), 
         .Z(n13128)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4586_3_lut.init = 16'hcaca;
    LUT4 i4585_3_lut (.A(\array[226] [1]), .B(\array[227] [1]), .C(r_addr[0]), 
         .Z(n13127)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4585_3_lut.init = 16'hcaca;
    LUT4 i4584_3_lut (.A(\array[224] [1]), .B(\array[225] [1]), .C(r_addr[0]), 
         .Z(n13126)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4584_3_lut.init = 16'hcaca;
    LUT4 i6349_3_lut (.A(\array[214] [0]), .B(\array[215] [0]), .C(r_addr[0]), 
         .Z(n14891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6349_3_lut.init = 16'hcaca;
    LUT4 i6348_3_lut (.A(\array[212] [0]), .B(\array[213] [0]), .C(r_addr[0]), 
         .Z(n14890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6348_3_lut.init = 16'hcaca;
    LUT4 i5495_3_lut (.A(\array[126] [5]), .B(\array[127] [5]), .C(r_addr[0]), 
         .Z(n14037)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5495_3_lut.init = 16'hcaca;
    LUT4 i5494_3_lut (.A(\array[124] [5]), .B(\array[125] [5]), .C(r_addr[0]), 
         .Z(n14036)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5494_3_lut.init = 16'hcaca;
    LUT4 i5493_3_lut (.A(\array[122] [5]), .B(\array[123] [5]), .C(r_addr[0]), 
         .Z(n14035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5493_3_lut.init = 16'hcaca;
    LUT4 i5492_3_lut (.A(\array[120] [5]), .B(\array[121] [5]), .C(r_addr[0]), 
         .Z(n14034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5492_3_lut.init = 16'hcaca;
    LUT4 i5491_3_lut (.A(\array[118] [5]), .B(\array[119] [5]), .C(r_addr[0]), 
         .Z(n14033)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5491_3_lut.init = 16'hcaca;
    LUT4 i5490_3_lut (.A(\array[116] [5]), .B(\array[117] [5]), .C(r_addr[0]), 
         .Z(n14032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5490_3_lut.init = 16'hcaca;
    LUT4 i5489_3_lut (.A(\array[114] [5]), .B(\array[115] [5]), .C(r_addr[0]), 
         .Z(n14031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5489_3_lut.init = 16'hcaca;
    LUT4 i5488_3_lut (.A(\array[112] [5]), .B(\array[113] [5]), .C(r_addr[0]), 
         .Z(n14030)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5488_3_lut.init = 16'hcaca;
    LUT4 i5487_3_lut (.A(\array[110] [5]), .B(\array[111] [5]), .C(r_addr[0]), 
         .Z(n14029)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5487_3_lut.init = 16'hcaca;
    LUT4 i5486_3_lut (.A(\array[108] [5]), .B(\array[109] [5]), .C(r_addr[0]), 
         .Z(n14028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5486_3_lut.init = 16'hcaca;
    LUT4 i5485_3_lut (.A(\array[106] [5]), .B(\array[107] [5]), .C(r_addr[0]), 
         .Z(n14027)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5485_3_lut.init = 16'hcaca;
    LUT4 i5484_3_lut (.A(\array[104] [5]), .B(\array[105] [5]), .C(r_addr[0]), 
         .Z(n14026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5484_3_lut.init = 16'hcaca;
    LUT4 i4568_3_lut (.A(\array[222] [1]), .B(\array[223] [1]), .C(r_addr[0]), 
         .Z(n13110)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4568_3_lut.init = 16'hcaca;
    LUT4 i4567_3_lut (.A(\array[220] [1]), .B(\array[221] [1]), .C(r_addr[0]), 
         .Z(n13109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4567_3_lut.init = 16'hcaca;
    LUT4 i5483_3_lut (.A(\array[102] [5]), .B(\array[103] [5]), .C(r_addr[0]), 
         .Z(n14025)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5483_3_lut.init = 16'hcaca;
    LUT4 i5482_3_lut (.A(\array[100] [5]), .B(\array[101] [5]), .C(r_addr[0]), 
         .Z(n14024)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5482_3_lut.init = 16'hcaca;
    LUT4 i4566_3_lut (.A(\array[218] [1]), .B(\array[219] [1]), .C(r_addr[0]), 
         .Z(n13108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4566_3_lut.init = 16'hcaca;
    LUT4 i4565_3_lut (.A(\array[216] [1]), .B(\array[217] [1]), .C(r_addr[0]), 
         .Z(n13107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4565_3_lut.init = 16'hcaca;
    LUT4 i4564_3_lut (.A(\array[214] [1]), .B(\array[215] [1]), .C(r_addr[0]), 
         .Z(n13106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4564_3_lut.init = 16'hcaca;
    LUT4 i4563_3_lut (.A(\array[212] [1]), .B(\array[213] [1]), .C(r_addr[0]), 
         .Z(n13105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4563_3_lut.init = 16'hcaca;
    LUT4 i5481_3_lut (.A(\array[98] [5]), .B(\array[99] [5]), .C(r_addr[0]), 
         .Z(n14023)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5481_3_lut.init = 16'hcaca;
    LUT4 i5480_3_lut (.A(\array[96] [5]), .B(\array[97] [5]), .C(r_addr[0]), 
         .Z(n14022)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5480_3_lut.init = 16'hcaca;
    LUT4 i4562_3_lut (.A(\array[210] [1]), .B(\array[211] [1]), .C(r_addr[0]), 
         .Z(n13104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4562_3_lut.init = 16'hcaca;
    LUT4 i4561_3_lut (.A(\array[208] [1]), .B(\array[209] [1]), .C(r_addr[0]), 
         .Z(n13103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4561_3_lut.init = 16'hcaca;
    LUT4 i4560_3_lut (.A(\array[206] [1]), .B(\array[207] [1]), .C(r_addr[0]), 
         .Z(n13102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4560_3_lut.init = 16'hcaca;
    LUT4 i4559_3_lut (.A(\array[204] [1]), .B(\array[205] [1]), .C(r_addr[0]), 
         .Z(n13101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4559_3_lut.init = 16'hcaca;
    LUT4 i4558_3_lut (.A(\array[202] [1]), .B(\array[203] [1]), .C(r_addr[0]), 
         .Z(n13100)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4558_3_lut.init = 16'hcaca;
    LUT4 i4557_3_lut (.A(\array[200] [1]), .B(\array[201] [1]), .C(r_addr[0]), 
         .Z(n13099)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4557_3_lut.init = 16'hcaca;
    LUT4 i4556_3_lut (.A(\array[198] [1]), .B(\array[199] [1]), .C(r_addr[0]), 
         .Z(n13098)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4556_3_lut.init = 16'hcaca;
    LUT4 i4555_3_lut (.A(\array[196] [1]), .B(\array[197] [1]), .C(r_addr[0]), 
         .Z(n13097)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4555_3_lut.init = 16'hcaca;
    LUT4 i4554_3_lut (.A(\array[194] [1]), .B(\array[195] [1]), .C(r_addr[0]), 
         .Z(n13096)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4554_3_lut.init = 16'hcaca;
    LUT4 i4553_3_lut (.A(\array[192] [1]), .B(\array[193] [1]), .C(r_addr[0]), 
         .Z(n13095)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4553_3_lut.init = 16'hcaca;
    LUT4 i6347_3_lut (.A(\array[210] [0]), .B(\array[211] [0]), .C(r_addr[0]), 
         .Z(n14889)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6347_3_lut.init = 16'hcaca;
    LUT4 i6346_3_lut (.A(\array[208] [0]), .B(\array[209] [0]), .C(r_addr[0]), 
         .Z(n14888)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6346_3_lut.init = 16'hcaca;
    LUT4 i6374_3_lut (.A(\array[234] [0]), .B(\array[235] [0]), .C(r_addr[0]), 
         .Z(n14916)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6374_3_lut.init = 16'hcaca;
    LUT4 i6373_3_lut (.A(\array[232] [0]), .B(\array[233] [0]), .C(r_addr[0]), 
         .Z(n14915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6373_3_lut.init = 16'hcaca;
    LUT4 i5943_3_lut (.A(\array[62] [7]), .B(\array[63] [7]), .C(r_addr[0]), 
         .Z(n14485)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5943_3_lut.init = 16'hcaca;
    LUT4 i5942_3_lut (.A(\array[60] [7]), .B(\array[61] [7]), .C(r_addr[0]), 
         .Z(n14484)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5942_3_lut.init = 16'hcaca;
    LUT4 i5941_3_lut (.A(\array[58] [7]), .B(\array[59] [7]), .C(r_addr[0]), 
         .Z(n14483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5941_3_lut.init = 16'hcaca;
    LUT4 i5940_3_lut (.A(\array[56] [7]), .B(\array[57] [7]), .C(r_addr[0]), 
         .Z(n14482)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5940_3_lut.init = 16'hcaca;
    LUT4 i5939_3_lut (.A(\array[54] [7]), .B(\array[55] [7]), .C(r_addr[0]), 
         .Z(n14481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5939_3_lut.init = 16'hcaca;
    LUT4 i5938_3_lut (.A(\array[52] [7]), .B(\array[53] [7]), .C(r_addr[0]), 
         .Z(n14480)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5938_3_lut.init = 16'hcaca;
    LUT4 i6291_3_lut (.A(\array[158] [0]), .B(\array[159] [0]), .C(r_addr[0]), 
         .Z(n14833)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6291_3_lut.init = 16'hcaca;
    LUT4 i6290_3_lut (.A(\array[156] [0]), .B(\array[157] [0]), .C(r_addr[0]), 
         .Z(n14832)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6290_3_lut.init = 16'hcaca;
    LUT4 i4537_3_lut (.A(\array[190] [1]), .B(\array[191] [1]), .C(r_addr[0]), 
         .Z(n13079)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4537_3_lut.init = 16'hcaca;
    LUT4 i4536_3_lut (.A(\array[188] [1]), .B(\array[189] [1]), .C(r_addr[0]), 
         .Z(n13078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4536_3_lut.init = 16'hcaca;
    LUT4 i4535_3_lut (.A(\array[186] [1]), .B(\array[187] [1]), .C(r_addr[0]), 
         .Z(n13077)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4535_3_lut.init = 16'hcaca;
    LUT4 i4534_3_lut (.A(\array[184] [1]), .B(\array[185] [1]), .C(r_addr[0]), 
         .Z(n13076)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4534_3_lut.init = 16'hcaca;
    LUT4 i5937_3_lut (.A(\array[50] [7]), .B(\array[51] [7]), .C(r_addr[0]), 
         .Z(n14479)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5937_3_lut.init = 16'hcaca;
    LUT4 i5936_3_lut (.A(\array[48] [7]), .B(\array[49] [7]), .C(r_addr[0]), 
         .Z(n14478)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5936_3_lut.init = 16'hcaca;
    LUT4 i4533_3_lut (.A(\array[182] [1]), .B(\array[183] [1]), .C(r_addr[0]), 
         .Z(n13075)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4533_3_lut.init = 16'hcaca;
    LUT4 i4532_3_lut (.A(\array[180] [1]), .B(\array[181] [1]), .C(r_addr[0]), 
         .Z(n13074)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4532_3_lut.init = 16'hcaca;
    LUT4 i4531_3_lut (.A(\array[178] [1]), .B(\array[179] [1]), .C(r_addr[0]), 
         .Z(n13073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4531_3_lut.init = 16'hcaca;
    LUT4 i4530_3_lut (.A(\array[176] [1]), .B(\array[177] [1]), .C(r_addr[0]), 
         .Z(n13072)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4530_3_lut.init = 16'hcaca;
    LUT4 i4529_3_lut (.A(\array[174] [1]), .B(\array[175] [1]), .C(r_addr[0]), 
         .Z(n13071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4529_3_lut.init = 16'hcaca;
    LUT4 i4528_3_lut (.A(\array[172] [1]), .B(\array[173] [1]), .C(r_addr[0]), 
         .Z(n13070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4528_3_lut.init = 16'hcaca;
    LUT4 i4527_3_lut (.A(\array[170] [1]), .B(\array[171] [1]), .C(r_addr[0]), 
         .Z(n13069)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4527_3_lut.init = 16'hcaca;
    LUT4 i4526_3_lut (.A(\array[168] [1]), .B(\array[169] [1]), .C(r_addr[0]), 
         .Z(n13068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4526_3_lut.init = 16'hcaca;
    LUT4 i5935_3_lut (.A(\array[46] [7]), .B(\array[47] [7]), .C(r_addr[0]), 
         .Z(n14477)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5935_3_lut.init = 16'hcaca;
    LUT4 i5934_3_lut (.A(\array[44] [7]), .B(\array[45] [7]), .C(r_addr[0]), 
         .Z(n14476)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5934_3_lut.init = 16'hcaca;
    LUT4 i4525_3_lut (.A(\array[166] [1]), .B(\array[167] [1]), .C(r_addr[0]), 
         .Z(n13067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4525_3_lut.init = 16'hcaca;
    LUT4 i4524_3_lut (.A(\array[164] [1]), .B(\array[165] [1]), .C(r_addr[0]), 
         .Z(n13066)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4524_3_lut.init = 16'hcaca;
    LUT4 i4523_3_lut (.A(\array[162] [1]), .B(\array[163] [1]), .C(r_addr[0]), 
         .Z(n13065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4523_3_lut.init = 16'hcaca;
    LUT4 i4522_3_lut (.A(\array[160] [1]), .B(\array[161] [1]), .C(r_addr[0]), 
         .Z(n13064)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4522_3_lut.init = 16'hcaca;
    LUT4 i5933_3_lut (.A(\array[42] [7]), .B(\array[43] [7]), .C(r_addr[0]), 
         .Z(n14475)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5933_3_lut.init = 16'hcaca;
    LUT4 i5932_3_lut (.A(\array[40] [7]), .B(\array[41] [7]), .C(r_addr[0]), 
         .Z(n14474)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5932_3_lut.init = 16'hcaca;
    LUT4 i5931_3_lut (.A(\array[38] [7]), .B(\array[39] [7]), .C(r_addr[0]), 
         .Z(n14473)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5931_3_lut.init = 16'hcaca;
    LUT4 i5930_3_lut (.A(\array[36] [7]), .B(\array[37] [7]), .C(r_addr[0]), 
         .Z(n14472)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5930_3_lut.init = 16'hcaca;
    LUT4 i6289_3_lut (.A(\array[154] [0]), .B(\array[155] [0]), .C(r_addr[0]), 
         .Z(n14831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6289_3_lut.init = 16'hcaca;
    LUT4 i6288_3_lut (.A(\array[152] [0]), .B(\array[153] [0]), .C(r_addr[0]), 
         .Z(n14830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6288_3_lut.init = 16'hcaca;
    LUT4 i6345_3_lut (.A(\array[206] [0]), .B(\array[207] [0]), .C(r_addr[0]), 
         .Z(n14887)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6345_3_lut.init = 16'hcaca;
    LUT4 i6344_3_lut (.A(\array[204] [0]), .B(\array[205] [0]), .C(r_addr[0]), 
         .Z(n14886)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6344_3_lut.init = 16'hcaca;
    LUT4 i5464_3_lut (.A(\array[94] [5]), .B(\array[95] [5]), .C(r_addr[0]), 
         .Z(n14006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5464_3_lut.init = 16'hcaca;
    LUT4 i5463_3_lut (.A(\array[92] [5]), .B(\array[93] [5]), .C(r_addr[0]), 
         .Z(n14005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5463_3_lut.init = 16'hcaca;
    LUT4 i5929_3_lut (.A(\array[34] [7]), .B(\array[35] [7]), .C(r_addr[0]), 
         .Z(n14471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5929_3_lut.init = 16'hcaca;
    LUT4 i5928_3_lut (.A(\array[32] [7]), .B(\array[33] [7]), .C(r_addr[0]), 
         .Z(n14470)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5928_3_lut.init = 16'hcaca;
    LUT4 i5462_3_lut (.A(\array[90] [5]), .B(\array[91] [5]), .C(r_addr[0]), 
         .Z(n14004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5462_3_lut.init = 16'hcaca;
    LUT4 i5461_3_lut (.A(\array[88] [5]), .B(\array[89] [5]), .C(r_addr[0]), 
         .Z(n14003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5461_3_lut.init = 16'hcaca;
    LUT4 i5460_3_lut (.A(\array[86] [5]), .B(\array[87] [5]), .C(r_addr[0]), 
         .Z(n14002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5460_3_lut.init = 16'hcaca;
    LUT4 i5459_3_lut (.A(\array[84] [5]), .B(\array[85] [5]), .C(r_addr[0]), 
         .Z(n14001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5459_3_lut.init = 16'hcaca;
    LUT4 i5458_3_lut (.A(\array[82] [5]), .B(\array[83] [5]), .C(r_addr[0]), 
         .Z(n14000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5458_3_lut.init = 16'hcaca;
    LUT4 i5457_3_lut (.A(\array[80] [5]), .B(\array[81] [5]), .C(r_addr[0]), 
         .Z(n13999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5457_3_lut.init = 16'hcaca;
    LUT4 i5456_3_lut (.A(\array[78] [5]), .B(\array[79] [5]), .C(r_addr[0]), 
         .Z(n13998)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5456_3_lut.init = 16'hcaca;
    LUT4 i5455_3_lut (.A(\array[76] [5]), .B(\array[77] [5]), .C(r_addr[0]), 
         .Z(n13997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5455_3_lut.init = 16'hcaca;
    LUT4 i5454_3_lut (.A(\array[74] [5]), .B(\array[75] [5]), .C(r_addr[0]), 
         .Z(n13996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5454_3_lut.init = 16'hcaca;
    LUT4 i5453_3_lut (.A(\array[72] [5]), .B(\array[73] [5]), .C(r_addr[0]), 
         .Z(n13995)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5453_3_lut.init = 16'hcaca;
    LUT4 i5452_3_lut (.A(\array[70] [5]), .B(\array[71] [5]), .C(r_addr[0]), 
         .Z(n13994)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5452_3_lut.init = 16'hcaca;
    LUT4 i5451_3_lut (.A(\array[68] [5]), .B(\array[69] [5]), .C(r_addr[0]), 
         .Z(n13993)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5451_3_lut.init = 16'hcaca;
    LUT4 i6287_3_lut (.A(\array[150] [0]), .B(\array[151] [0]), .C(r_addr[0]), 
         .Z(n14829)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6287_3_lut.init = 16'hcaca;
    LUT4 i6286_3_lut (.A(\array[148] [0]), .B(\array[149] [0]), .C(r_addr[0]), 
         .Z(n14828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6286_3_lut.init = 16'hcaca;
    LUT4 i5450_3_lut (.A(\array[66] [5]), .B(\array[67] [5]), .C(r_addr[0]), 
         .Z(n13992)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5450_3_lut.init = 16'hcaca;
    LUT4 i5449_3_lut (.A(\array[64] [5]), .B(\array[65] [5]), .C(r_addr[0]), 
         .Z(n13991)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5449_3_lut.init = 16'hcaca;
    LUT4 i6285_3_lut (.A(\array[146] [0]), .B(\array[147] [0]), .C(r_addr[0]), 
         .Z(n14827)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6285_3_lut.init = 16'hcaca;
    LUT4 i6284_3_lut (.A(\array[144] [0]), .B(\array[145] [0]), .C(r_addr[0]), 
         .Z(n14826)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6284_3_lut.init = 16'hcaca;
    LUT4 i6343_3_lut (.A(\array[202] [0]), .B(\array[203] [0]), .C(r_addr[0]), 
         .Z(n14885)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6343_3_lut.init = 16'hcaca;
    LUT4 i6342_3_lut (.A(\array[200] [0]), .B(\array[201] [0]), .C(r_addr[0]), 
         .Z(n14884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6342_3_lut.init = 16'hcaca;
    LUT4 i6372_3_lut (.A(\array[230] [0]), .B(\array[231] [0]), .C(r_addr[0]), 
         .Z(n14914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6372_3_lut.init = 16'hcaca;
    LUT4 i6371_3_lut (.A(\array[228] [0]), .B(\array[229] [0]), .C(r_addr[0]), 
         .Z(n14913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6371_3_lut.init = 16'hcaca;
    LUT4 i6167_3_lut (.A(\array[30] [0]), .B(\array[31] [0]), .C(r_addr[0]), 
         .Z(n14709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6167_3_lut.init = 16'hcaca;
    LUT4 i6166_3_lut (.A(\array[28] [0]), .B(\array[29] [0]), .C(r_addr[0]), 
         .Z(n14708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6166_3_lut.init = 16'hcaca;
    LUT4 i6165_3_lut (.A(\array[26] [0]), .B(\array[27] [0]), .C(r_addr[0]), 
         .Z(n14707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6165_3_lut.init = 16'hcaca;
    LUT4 i6164_3_lut (.A(\array[24] [0]), .B(\array[25] [0]), .C(r_addr[0]), 
         .Z(n14706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6164_3_lut.init = 16'hcaca;
    LUT4 i6283_3_lut (.A(\array[142] [0]), .B(\array[143] [0]), .C(r_addr[0]), 
         .Z(n14825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6283_3_lut.init = 16'hcaca;
    LUT4 i6282_3_lut (.A(\array[140] [0]), .B(\array[141] [0]), .C(r_addr[0]), 
         .Z(n14824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6282_3_lut.init = 16'hcaca;
    LUT4 i6163_3_lut (.A(\array[22] [0]), .B(\array[23] [0]), .C(r_addr[0]), 
         .Z(n14705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6163_3_lut.init = 16'hcaca;
    LUT4 i6162_3_lut (.A(\array[20] [0]), .B(\array[21] [0]), .C(r_addr[0]), 
         .Z(n14704)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6162_3_lut.init = 16'hcaca;
    LUT4 i5433_3_lut (.A(\array[62] [5]), .B(\array[63] [5]), .C(r_addr[0]), 
         .Z(n13975)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5433_3_lut.init = 16'hcaca;
    LUT4 i5432_3_lut (.A(\array[60] [5]), .B(\array[61] [5]), .C(r_addr[0]), 
         .Z(n13974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5432_3_lut.init = 16'hcaca;
    LUT4 i6161_3_lut (.A(\array[18] [0]), .B(\array[19] [0]), .C(r_addr[0]), 
         .Z(n14703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6161_3_lut.init = 16'hcaca;
    LUT4 i6160_3_lut (.A(\array[16] [0]), .B(\array[17] [0]), .C(r_addr[0]), 
         .Z(n14702)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6160_3_lut.init = 16'hcaca;
    LUT4 i6281_3_lut (.A(\array[138] [0]), .B(\array[139] [0]), .C(r_addr[0]), 
         .Z(n14823)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6281_3_lut.init = 16'hcaca;
    LUT4 i6280_3_lut (.A(\array[136] [0]), .B(\array[137] [0]), .C(r_addr[0]), 
         .Z(n14822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6280_3_lut.init = 16'hcaca;
    LUT4 i6341_3_lut (.A(\array[198] [0]), .B(\array[199] [0]), .C(r_addr[0]), 
         .Z(n14883)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6341_3_lut.init = 16'hcaca;
    LUT4 i6340_3_lut (.A(\array[196] [0]), .B(\array[197] [0]), .C(r_addr[0]), 
         .Z(n14882)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6340_3_lut.init = 16'hcaca;
    LUT4 i5431_3_lut (.A(\array[58] [5]), .B(\array[59] [5]), .C(r_addr[0]), 
         .Z(n13973)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5431_3_lut.init = 16'hcaca;
    LUT4 i5430_3_lut (.A(\array[56] [5]), .B(\array[57] [5]), .C(r_addr[0]), 
         .Z(n13972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5430_3_lut.init = 16'hcaca;
    LUT4 i5429_3_lut (.A(\array[54] [5]), .B(\array[55] [5]), .C(r_addr[0]), 
         .Z(n13971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5429_3_lut.init = 16'hcaca;
    LUT4 i5428_3_lut (.A(\array[52] [5]), .B(\array[53] [5]), .C(r_addr[0]), 
         .Z(n13970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5428_3_lut.init = 16'hcaca;
    LUT4 i5427_3_lut (.A(\array[50] [5]), .B(\array[51] [5]), .C(r_addr[0]), 
         .Z(n13969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5427_3_lut.init = 16'hcaca;
    LUT4 i5426_3_lut (.A(\array[48] [5]), .B(\array[49] [5]), .C(r_addr[0]), 
         .Z(n13968)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5426_3_lut.init = 16'hcaca;
    LUT4 i5425_3_lut (.A(\array[46] [5]), .B(\array[47] [5]), .C(r_addr[0]), 
         .Z(n13967)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5425_3_lut.init = 16'hcaca;
    LUT4 i5424_3_lut (.A(\array[44] [5]), .B(\array[45] [5]), .C(r_addr[0]), 
         .Z(n13966)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5424_3_lut.init = 16'hcaca;
    LUT4 i6159_3_lut (.A(\array[14] [0]), .B(\array[15] [0]), .C(r_addr[0]), 
         .Z(n14701)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6159_3_lut.init = 16'hcaca;
    LUT4 i6158_3_lut (.A(\array[12] [0]), .B(\array[13] [0]), .C(r_addr[0]), 
         .Z(n14700)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6158_3_lut.init = 16'hcaca;
    LUT4 i5423_3_lut (.A(\array[42] [5]), .B(\array[43] [5]), .C(r_addr[0]), 
         .Z(n13965)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5423_3_lut.init = 16'hcaca;
    LUT4 i5422_3_lut (.A(\array[40] [5]), .B(\array[41] [5]), .C(r_addr[0]), 
         .Z(n13964)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5422_3_lut.init = 16'hcaca;
    LUT4 i5421_3_lut (.A(\array[38] [5]), .B(\array[39] [5]), .C(r_addr[0]), 
         .Z(n13963)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5421_3_lut.init = 16'hcaca;
    LUT4 i5420_3_lut (.A(\array[36] [5]), .B(\array[37] [5]), .C(r_addr[0]), 
         .Z(n13962)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5420_3_lut.init = 16'hcaca;
    LUT4 i5419_3_lut (.A(\array[34] [5]), .B(\array[35] [5]), .C(r_addr[0]), 
         .Z(n13961)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5419_3_lut.init = 16'hcaca;
    LUT4 i5418_3_lut (.A(\array[32] [5]), .B(\array[33] [5]), .C(r_addr[0]), 
         .Z(n13960)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5418_3_lut.init = 16'hcaca;
    LUT4 i6157_3_lut (.A(\array[10] [0]), .B(\array[11] [0]), .C(r_addr[0]), 
         .Z(n14699)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6157_3_lut.init = 16'hcaca;
    LUT4 i6156_3_lut (.A(\array[8] [0]), .B(\array[9] [0]), .C(r_addr[0]), 
         .Z(n14698)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6156_3_lut.init = 16'hcaca;
    LUT4 i6279_3_lut (.A(\array[134] [0]), .B(\array[135] [0]), .C(r_addr[0]), 
         .Z(n14821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6279_3_lut.init = 16'hcaca;
    LUT4 i6278_3_lut (.A(\array[132] [0]), .B(\array[133] [0]), .C(r_addr[0]), 
         .Z(n14820)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6278_3_lut.init = 16'hcaca;
    LUT4 i6155_3_lut (.A(\array[6] [0]), .B(\array[7] [0]), .C(r_addr[0]), 
         .Z(n14697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6155_3_lut.init = 16'hcaca;
    LUT4 i6154_3_lut (.A(\array[4] [0]), .B(\array[5] [0]), .C(r_addr[0]), 
         .Z(n14696)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6154_3_lut.init = 16'hcaca;
    LUT4 i4506_3_lut (.A(\array[158] [1]), .B(\array[159] [1]), .C(r_addr[0]), 
         .Z(n13048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4506_3_lut.init = 16'hcaca;
    LUT4 i4505_3_lut (.A(\array[156] [1]), .B(\array[157] [1]), .C(r_addr[0]), 
         .Z(n13047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4505_3_lut.init = 16'hcaca;
    LUT4 i4504_3_lut (.A(\array[154] [1]), .B(\array[155] [1]), .C(r_addr[0]), 
         .Z(n13046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4504_3_lut.init = 16'hcaca;
    LUT4 i4503_3_lut (.A(\array[152] [1]), .B(\array[153] [1]), .C(r_addr[0]), 
         .Z(n13045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4503_3_lut.init = 16'hcaca;
    LUT4 i4502_3_lut (.A(\array[150] [1]), .B(\array[151] [1]), .C(r_addr[0]), 
         .Z(n13044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4502_3_lut.init = 16'hcaca;
    LUT4 i4501_3_lut (.A(\array[148] [1]), .B(\array[149] [1]), .C(r_addr[0]), 
         .Z(n13043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4501_3_lut.init = 16'hcaca;
    LUT4 i4500_3_lut (.A(\array[146] [1]), .B(\array[147] [1]), .C(r_addr[0]), 
         .Z(n13042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4500_3_lut.init = 16'hcaca;
    LUT4 i4499_3_lut (.A(\array[144] [1]), .B(\array[145] [1]), .C(r_addr[0]), 
         .Z(n13041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4499_3_lut.init = 16'hcaca;
    LUT4 i4498_3_lut (.A(\array[142] [1]), .B(\array[143] [1]), .C(r_addr[0]), 
         .Z(n13040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4498_3_lut.init = 16'hcaca;
    LUT4 i4497_3_lut (.A(\array[140] [1]), .B(\array[141] [1]), .C(r_addr[0]), 
         .Z(n13039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4497_3_lut.init = 16'hcaca;
    LUT4 i4496_3_lut (.A(\array[138] [1]), .B(\array[139] [1]), .C(r_addr[0]), 
         .Z(n13038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4496_3_lut.init = 16'hcaca;
    LUT4 i4495_3_lut (.A(\array[136] [1]), .B(\array[137] [1]), .C(r_addr[0]), 
         .Z(n13037)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4495_3_lut.init = 16'hcaca;
    LUT4 i4494_3_lut (.A(\array[134] [1]), .B(\array[135] [1]), .C(r_addr[0]), 
         .Z(n13036)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4494_3_lut.init = 16'hcaca;
    LUT4 i4493_3_lut (.A(\array[132] [1]), .B(\array[133] [1]), .C(r_addr[0]), 
         .Z(n13035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4493_3_lut.init = 16'hcaca;
    LUT4 i4492_3_lut (.A(\array[130] [1]), .B(\array[131] [1]), .C(r_addr[0]), 
         .Z(n13034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4492_3_lut.init = 16'hcaca;
    LUT4 i4491_3_lut (.A(\array[128] [1]), .B(\array[129] [1]), .C(r_addr[0]), 
         .Z(n13033)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4491_3_lut.init = 16'hcaca;
    LUT4 i5912_3_lut (.A(\array[30] [7]), .B(\array[31] [7]), .C(r_addr[0]), 
         .Z(n14454)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5912_3_lut.init = 16'hcaca;
    LUT4 i5911_3_lut (.A(\array[28] [7]), .B(\array[29] [7]), .C(r_addr[0]), 
         .Z(n14453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5911_3_lut.init = 16'hcaca;
    LUT4 i6153_3_lut (.A(\array[2] [0]), .B(\array[3] [0]), .C(r_addr[0]), 
         .Z(n14695)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6153_3_lut.init = 16'hcaca;
    LUT4 i6152_3_lut (.A(\array[0] [0]), .B(\array[1] [0]), .C(r_addr[0]), 
         .Z(n14694)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6152_3_lut.init = 16'hcaca;
    LUT4 i6277_3_lut (.A(\array[130] [0]), .B(\array[131] [0]), .C(r_addr[0]), 
         .Z(n14819)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6277_3_lut.init = 16'hcaca;
    LUT4 i6276_3_lut (.A(\array[128] [0]), .B(\array[129] [0]), .C(r_addr[0]), 
         .Z(n14818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6276_3_lut.init = 16'hcaca;
    LUT4 i6339_3_lut (.A(\array[194] [0]), .B(\array[195] [0]), .C(r_addr[0]), 
         .Z(n14881)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6339_3_lut.init = 16'hcaca;
    LUT4 i6338_3_lut (.A(\array[192] [0]), .B(\array[193] [0]), .C(r_addr[0]), 
         .Z(n14880)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6338_3_lut.init = 16'hcaca;
    LUT4 i6370_3_lut (.A(\array[226] [0]), .B(\array[227] [0]), .C(r_addr[0]), 
         .Z(n14912)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6370_3_lut.init = 16'hcaca;
    LUT4 i6369_3_lut (.A(\array[224] [0]), .B(\array[225] [0]), .C(r_addr[0]), 
         .Z(n14911)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6369_3_lut.init = 16'hcaca;
    LUT4 i5910_3_lut (.A(\array[26] [7]), .B(\array[27] [7]), .C(r_addr[0]), 
         .Z(n14452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5910_3_lut.init = 16'hcaca;
    LUT4 i5909_3_lut (.A(\array[24] [7]), .B(\array[25] [7]), .C(r_addr[0]), 
         .Z(n14451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5909_3_lut.init = 16'hcaca;
    LUT4 i5908_3_lut (.A(\array[22] [7]), .B(\array[23] [7]), .C(r_addr[0]), 
         .Z(n14450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5908_3_lut.init = 16'hcaca;
    LUT4 i5907_3_lut (.A(\array[20] [7]), .B(\array[21] [7]), .C(r_addr[0]), 
         .Z(n14449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5907_3_lut.init = 16'hcaca;
    LUT4 i5906_3_lut (.A(\array[18] [7]), .B(\array[19] [7]), .C(r_addr[0]), 
         .Z(n14448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5906_3_lut.init = 16'hcaca;
    LUT4 i5905_3_lut (.A(\array[16] [7]), .B(\array[17] [7]), .C(r_addr[0]), 
         .Z(n14447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5905_3_lut.init = 16'hcaca;
    LUT4 i5904_3_lut (.A(\array[14] [7]), .B(\array[15] [7]), .C(r_addr[0]), 
         .Z(n14446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5904_3_lut.init = 16'hcaca;
    LUT4 i5903_3_lut (.A(\array[12] [7]), .B(\array[13] [7]), .C(r_addr[0]), 
         .Z(n14445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5903_3_lut.init = 16'hcaca;
    LUT4 i5902_3_lut (.A(\array[10] [7]), .B(\array[11] [7]), .C(r_addr[0]), 
         .Z(n14444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5902_3_lut.init = 16'hcaca;
    LUT4 i5901_3_lut (.A(\array[8] [7]), .B(\array[9] [7]), .C(r_addr[0]), 
         .Z(n14443)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5901_3_lut.init = 16'hcaca;
    LUT4 i4475_3_lut (.A(\array[126] [1]), .B(\array[127] [1]), .C(r_addr[0]), 
         .Z(n13017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4475_3_lut.init = 16'hcaca;
    LUT4 i4474_3_lut (.A(\array[124] [1]), .B(\array[125] [1]), .C(r_addr[0]), 
         .Z(n13016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4474_3_lut.init = 16'hcaca;
    LUT4 i5900_3_lut (.A(\array[6] [7]), .B(\array[7] [7]), .C(r_addr[0]), 
         .Z(n14442)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5900_3_lut.init = 16'hcaca;
    LUT4 i5899_3_lut (.A(\array[4] [7]), .B(\array[5] [7]), .C(r_addr[0]), 
         .Z(n14441)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5899_3_lut.init = 16'hcaca;
    LUT4 i4473_3_lut (.A(\array[122] [1]), .B(\array[123] [1]), .C(r_addr[0]), 
         .Z(n13015)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4473_3_lut.init = 16'hcaca;
    LUT4 i4472_3_lut (.A(\array[120] [1]), .B(\array[121] [1]), .C(r_addr[0]), 
         .Z(n13014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4472_3_lut.init = 16'hcaca;
    LUT4 i4471_3_lut (.A(\array[118] [1]), .B(\array[119] [1]), .C(r_addr[0]), 
         .Z(n13013)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4471_3_lut.init = 16'hcaca;
    LUT4 i4470_3_lut (.A(\array[116] [1]), .B(\array[117] [1]), .C(r_addr[0]), 
         .Z(n13012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4470_3_lut.init = 16'hcaca;
    LUT4 i4469_3_lut (.A(\array[114] [1]), .B(\array[115] [1]), .C(r_addr[0]), 
         .Z(n13011)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4469_3_lut.init = 16'hcaca;
    LUT4 i4468_3_lut (.A(\array[112] [1]), .B(\array[113] [1]), .C(r_addr[0]), 
         .Z(n13010)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4468_3_lut.init = 16'hcaca;
    LUT4 i4467_3_lut (.A(\array[110] [1]), .B(\array[111] [1]), .C(r_addr[0]), 
         .Z(n13009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4467_3_lut.init = 16'hcaca;
    LUT4 i4466_3_lut (.A(\array[108] [1]), .B(\array[109] [1]), .C(r_addr[0]), 
         .Z(n13008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4466_3_lut.init = 16'hcaca;
    LUT4 i5402_3_lut (.A(\array[30] [5]), .B(\array[31] [5]), .C(r_addr[0]), 
         .Z(n13944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5402_3_lut.init = 16'hcaca;
    LUT4 i5401_3_lut (.A(\array[28] [5]), .B(\array[29] [5]), .C(r_addr[0]), 
         .Z(n13943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5401_3_lut.init = 16'hcaca;
    LUT4 i5898_3_lut (.A(\array[2] [7]), .B(\array[3] [7]), .C(r_addr[0]), 
         .Z(n14440)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5898_3_lut.init = 16'hcaca;
    LUT4 i5897_3_lut (.A(\array[0] [7]), .B(\array[1] [7]), .C(r_addr[0]), 
         .Z(n14439)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5897_3_lut.init = 16'hcaca;
    LUT4 i4465_3_lut (.A(\array[106] [1]), .B(\array[107] [1]), .C(r_addr[0]), 
         .Z(n13007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4465_3_lut.init = 16'hcaca;
    LUT4 i4464_3_lut (.A(\array[104] [1]), .B(\array[105] [1]), .C(r_addr[0]), 
         .Z(n13006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4464_3_lut.init = 16'hcaca;
    LUT4 i4463_3_lut (.A(\array[102] [1]), .B(\array[103] [1]), .C(r_addr[0]), 
         .Z(n13005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4463_3_lut.init = 16'hcaca;
    LUT4 i4462_3_lut (.A(\array[100] [1]), .B(\array[101] [1]), .C(r_addr[0]), 
         .Z(n13004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4462_3_lut.init = 16'hcaca;
    LUT4 i5400_3_lut (.A(\array[26] [5]), .B(\array[27] [5]), .C(r_addr[0]), 
         .Z(n13942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5400_3_lut.init = 16'hcaca;
    LUT4 i5399_3_lut (.A(\array[24] [5]), .B(\array[25] [5]), .C(r_addr[0]), 
         .Z(n13941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5399_3_lut.init = 16'hcaca;
    LUT4 i4461_3_lut (.A(\array[98] [1]), .B(\array[99] [1]), .C(r_addr[0]), 
         .Z(n13003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4461_3_lut.init = 16'hcaca;
    LUT4 i4460_3_lut (.A(\array[96] [1]), .B(\array[97] [1]), .C(r_addr[0]), 
         .Z(n13002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4460_3_lut.init = 16'hcaca;
    LUT4 i5398_3_lut (.A(\array[22] [5]), .B(\array[23] [5]), .C(r_addr[0]), 
         .Z(n13940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5398_3_lut.init = 16'hcaca;
    LUT4 i5397_3_lut (.A(\array[20] [5]), .B(\array[21] [5]), .C(r_addr[0]), 
         .Z(n13939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5397_3_lut.init = 16'hcaca;
    LUT4 i5396_3_lut (.A(\array[18] [5]), .B(\array[19] [5]), .C(r_addr[0]), 
         .Z(n13938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5396_3_lut.init = 16'hcaca;
    LUT4 i5395_3_lut (.A(\array[16] [5]), .B(\array[17] [5]), .C(r_addr[0]), 
         .Z(n13937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5395_3_lut.init = 16'hcaca;
    LUT4 i5394_3_lut (.A(\array[14] [5]), .B(\array[15] [5]), .C(r_addr[0]), 
         .Z(n13936)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5394_3_lut.init = 16'hcaca;
    LUT4 i5393_3_lut (.A(\array[12] [5]), .B(\array[13] [5]), .C(r_addr[0]), 
         .Z(n13935)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5393_3_lut.init = 16'hcaca;
    LUT4 i5392_3_lut (.A(\array[10] [5]), .B(\array[11] [5]), .C(r_addr[0]), 
         .Z(n13934)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5392_3_lut.init = 16'hcaca;
    LUT4 i5391_3_lut (.A(\array[8] [5]), .B(\array[9] [5]), .C(r_addr[0]), 
         .Z(n13933)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5391_3_lut.init = 16'hcaca;
    LUT4 i5390_3_lut (.A(\array[6] [5]), .B(\array[7] [5]), .C(r_addr[0]), 
         .Z(n13932)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5390_3_lut.init = 16'hcaca;
    LUT4 i5389_3_lut (.A(\array[4] [5]), .B(\array[5] [5]), .C(r_addr[0]), 
         .Z(n13931)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5389_3_lut.init = 16'hcaca;
    LUT4 i5388_3_lut (.A(\array[2] [5]), .B(\array[3] [5]), .C(r_addr[0]), 
         .Z(n13930)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5388_3_lut.init = 16'hcaca;
    LUT4 i5387_3_lut (.A(\array[0] [5]), .B(\array[1] [5]), .C(r_addr[0]), 
         .Z(n13929)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5387_3_lut.init = 16'hcaca;
    LUT4 i4444_3_lut (.A(\array[94] [1]), .B(\array[95] [1]), .C(r_addr[0]), 
         .Z(n12986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4444_3_lut.init = 16'hcaca;
    LUT4 i4443_3_lut (.A(\array[92] [1]), .B(\array[93] [1]), .C(r_addr[0]), 
         .Z(n12985)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4443_3_lut.init = 16'hcaca;
    LUT4 i4442_3_lut (.A(\array[90] [1]), .B(\array[91] [1]), .C(r_addr[0]), 
         .Z(n12984)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4442_3_lut.init = 16'hcaca;
    LUT4 i4441_3_lut (.A(\array[88] [1]), .B(\array[89] [1]), .C(r_addr[0]), 
         .Z(n12983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4441_3_lut.init = 16'hcaca;
    LUT4 i4440_3_lut (.A(\array[86] [1]), .B(\array[87] [1]), .C(r_addr[0]), 
         .Z(n12982)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4440_3_lut.init = 16'hcaca;
    LUT4 i4439_3_lut (.A(\array[84] [1]), .B(\array[85] [1]), .C(r_addr[0]), 
         .Z(n12981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4439_3_lut.init = 16'hcaca;
    LUT4 i4438_3_lut (.A(\array[82] [1]), .B(\array[83] [1]), .C(r_addr[0]), 
         .Z(n12980)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4438_3_lut.init = 16'hcaca;
    LUT4 i4437_3_lut (.A(\array[80] [1]), .B(\array[81] [1]), .C(r_addr[0]), 
         .Z(n12979)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4437_3_lut.init = 16'hcaca;
    LUT4 i4436_3_lut (.A(\array[78] [1]), .B(\array[79] [1]), .C(r_addr[0]), 
         .Z(n12978)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4436_3_lut.init = 16'hcaca;
    LUT4 i4435_3_lut (.A(\array[76] [1]), .B(\array[77] [1]), .C(r_addr[0]), 
         .Z(n12977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4435_3_lut.init = 16'hcaca;
    LUT4 i4434_3_lut (.A(\array[74] [1]), .B(\array[75] [1]), .C(r_addr[0]), 
         .Z(n12976)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4434_3_lut.init = 16'hcaca;
    LUT4 i4433_3_lut (.A(\array[72] [1]), .B(\array[73] [1]), .C(r_addr[0]), 
         .Z(n12975)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4433_3_lut.init = 16'hcaca;
    LUT4 i4432_3_lut (.A(\array[70] [1]), .B(\array[71] [1]), .C(r_addr[0]), 
         .Z(n12974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4432_3_lut.init = 16'hcaca;
    LUT4 i4431_3_lut (.A(\array[68] [1]), .B(\array[69] [1]), .C(r_addr[0]), 
         .Z(n12973)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4431_3_lut.init = 16'hcaca;
    LUT4 i4430_3_lut (.A(\array[66] [1]), .B(\array[67] [1]), .C(r_addr[0]), 
         .Z(n12972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4430_3_lut.init = 16'hcaca;
    LUT4 i4429_3_lut (.A(\array[64] [1]), .B(\array[65] [1]), .C(r_addr[0]), 
         .Z(n12971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4429_3_lut.init = 16'hcaca;
    LUT4 i4413_3_lut (.A(\array[62] [1]), .B(\array[63] [1]), .C(r_addr[0]), 
         .Z(n12955)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4413_3_lut.init = 16'hcaca;
    LUT4 i4412_3_lut (.A(\array[60] [1]), .B(\array[61] [1]), .C(r_addr[0]), 
         .Z(n12954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4412_3_lut.init = 16'hcaca;
    LUT4 i4411_3_lut (.A(\array[58] [1]), .B(\array[59] [1]), .C(r_addr[0]), 
         .Z(n12953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4411_3_lut.init = 16'hcaca;
    LUT4 i4410_3_lut (.A(\array[56] [1]), .B(\array[57] [1]), .C(r_addr[0]), 
         .Z(n12952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4410_3_lut.init = 16'hcaca;
    LUT4 i4409_3_lut (.A(\array[54] [1]), .B(\array[55] [1]), .C(r_addr[0]), 
         .Z(n12951)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4409_3_lut.init = 16'hcaca;
    LUT4 i4408_3_lut (.A(\array[52] [1]), .B(\array[53] [1]), .C(r_addr[0]), 
         .Z(n12950)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4408_3_lut.init = 16'hcaca;
    LUT4 i4407_3_lut (.A(\array[50] [1]), .B(\array[51] [1]), .C(r_addr[0]), 
         .Z(n12949)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4407_3_lut.init = 16'hcaca;
    LUT4 i4406_3_lut (.A(\array[48] [1]), .B(\array[49] [1]), .C(r_addr[0]), 
         .Z(n12948)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4406_3_lut.init = 16'hcaca;
    LUT4 i4405_3_lut (.A(\array[46] [1]), .B(\array[47] [1]), .C(r_addr[0]), 
         .Z(n12947)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4405_3_lut.init = 16'hcaca;
    LUT4 i4404_3_lut (.A(\array[44] [1]), .B(\array[45] [1]), .C(r_addr[0]), 
         .Z(n12946)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4404_3_lut.init = 16'hcaca;
    LUT4 i4403_3_lut (.A(\array[42] [1]), .B(\array[43] [1]), .C(r_addr[0]), 
         .Z(n12945)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4403_3_lut.init = 16'hcaca;
    LUT4 i4402_3_lut (.A(\array[40] [1]), .B(\array[41] [1]), .C(r_addr[0]), 
         .Z(n12944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4402_3_lut.init = 16'hcaca;
    LUT4 i4401_3_lut (.A(\array[38] [1]), .B(\array[39] [1]), .C(r_addr[0]), 
         .Z(n12943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4401_3_lut.init = 16'hcaca;
    LUT4 i4400_3_lut (.A(\array[36] [1]), .B(\array[37] [1]), .C(r_addr[0]), 
         .Z(n12942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4400_3_lut.init = 16'hcaca;
    LUT4 i4399_3_lut (.A(\array[34] [1]), .B(\array[35] [1]), .C(r_addr[0]), 
         .Z(n12941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4399_3_lut.init = 16'hcaca;
    LUT4 i4398_3_lut (.A(\array[32] [1]), .B(\array[33] [1]), .C(r_addr[0]), 
         .Z(n12940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4398_3_lut.init = 16'hcaca;
    LUT4 i5364_3_lut (.A(\array[254] [4]), .B(\array[255] [4]), .C(r_addr[0]), 
         .Z(n13906)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5364_3_lut.init = 16'hcaca;
    LUT4 i5363_3_lut (.A(\array[252] [4]), .B(\array[253] [4]), .C(r_addr[0]), 
         .Z(n13905)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5363_3_lut.init = 16'hcaca;
    LUT4 i5362_3_lut (.A(\array[250] [4]), .B(\array[251] [4]), .C(r_addr[0]), 
         .Z(n13904)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5362_3_lut.init = 16'hcaca;
    LUT4 i5361_3_lut (.A(\array[248] [4]), .B(\array[249] [4]), .C(r_addr[0]), 
         .Z(n13903)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5361_3_lut.init = 16'hcaca;
    LUT4 i5360_3_lut (.A(\array[246] [4]), .B(\array[247] [4]), .C(r_addr[0]), 
         .Z(n13902)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5360_3_lut.init = 16'hcaca;
    LUT4 i5359_3_lut (.A(\array[244] [4]), .B(\array[245] [4]), .C(r_addr[0]), 
         .Z(n13901)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5359_3_lut.init = 16'hcaca;
    LUT4 i5358_3_lut (.A(\array[242] [4]), .B(\array[243] [4]), .C(r_addr[0]), 
         .Z(n13900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5358_3_lut.init = 16'hcaca;
    LUT4 i5357_3_lut (.A(\array[240] [4]), .B(\array[241] [4]), .C(r_addr[0]), 
         .Z(n13899)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5357_3_lut.init = 16'hcaca;
    LUT4 i5356_3_lut (.A(\array[238] [4]), .B(\array[239] [4]), .C(maxfan_replicated_net_23), 
         .Z(n13898)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5356_3_lut.init = 16'hcaca;
    LUT4 i5355_3_lut (.A(\array[236] [4]), .B(\array[237] [4]), .C(maxfan_replicated_net_23), 
         .Z(n13897)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5355_3_lut.init = 16'hcaca;
    LUT4 i5354_3_lut (.A(\array[234] [4]), .B(\array[235] [4]), .C(maxfan_replicated_net_23), 
         .Z(n13896)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5354_3_lut.init = 16'hcaca;
    LUT4 i5353_3_lut (.A(\array[232] [4]), .B(\array[233] [4]), .C(maxfan_replicated_net_23), 
         .Z(n13895)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5353_3_lut.init = 16'hcaca;
    LUT4 i4382_3_lut (.A(\array[30] [1]), .B(\array[31] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4382_3_lut.init = 16'hcaca;
    LUT4 i4381_3_lut (.A(\array[28] [1]), .B(\array[29] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4381_3_lut.init = 16'hcaca;
    LUT4 i5352_3_lut (.A(\array[230] [4]), .B(\array[231] [4]), .C(maxfan_replicated_net_23), 
         .Z(n13894)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5352_3_lut.init = 16'hcaca;
    LUT4 i5351_3_lut (.A(\array[228] [4]), .B(\array[229] [4]), .C(maxfan_replicated_net_23), 
         .Z(n13893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5351_3_lut.init = 16'hcaca;
    LUT4 i4380_3_lut (.A(\array[26] [1]), .B(\array[27] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4380_3_lut.init = 16'hcaca;
    LUT4 i4379_3_lut (.A(\array[24] [1]), .B(\array[25] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12921)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4379_3_lut.init = 16'hcaca;
    LUT4 i4378_3_lut (.A(\array[22] [1]), .B(\array[23] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4378_3_lut.init = 16'hcaca;
    LUT4 i4377_3_lut (.A(\array[20] [1]), .B(\array[21] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12919)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4377_3_lut.init = 16'hcaca;
    LUT4 i5350_3_lut (.A(\array[226] [4]), .B(\array[227] [4]), .C(maxfan_replicated_net_23), 
         .Z(n13892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5350_3_lut.init = 16'hcaca;
    LUT4 i5349_3_lut (.A(\array[224] [4]), .B(\array[225] [4]), .C(maxfan_replicated_net_23), 
         .Z(n13891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5349_3_lut.init = 16'hcaca;
    LUT4 i4376_3_lut (.A(\array[18] [1]), .B(\array[19] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12918)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4376_3_lut.init = 16'hcaca;
    LUT4 i4375_3_lut (.A(\array[16] [1]), .B(\array[17] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12917)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4375_3_lut.init = 16'hcaca;
    LUT4 i4374_3_lut (.A(\array[14] [1]), .B(\array[15] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12916)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4374_3_lut.init = 16'hcaca;
    LUT4 i4373_3_lut (.A(\array[12] [1]), .B(\array[13] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4373_3_lut.init = 16'hcaca;
    LUT4 i4372_3_lut (.A(\array[10] [1]), .B(\array[11] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4372_3_lut.init = 16'hcaca;
    LUT4 i4371_3_lut (.A(\array[8] [1]), .B(\array[9] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4371_3_lut.init = 16'hcaca;
    LUT4 i4370_3_lut (.A(\array[6] [1]), .B(\array[7] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12912)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4370_3_lut.init = 16'hcaca;
    LUT4 i4369_3_lut (.A(\array[4] [1]), .B(\array[5] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12911)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4369_3_lut.init = 16'hcaca;
    LUT4 i4368_3_lut (.A(\array[2] [1]), .B(\array[3] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12910)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4368_3_lut.init = 16'hcaca;
    LUT4 i4367_3_lut (.A(\array[0] [1]), .B(\array[1] [1]), .C(maxfan_replicated_net_23), 
         .Z(n12909)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4367_3_lut.init = 16'hcaca;
    LUT4 i6144_3_lut (.A(n14684), .B(n14685), .C(r_addr[4]), .Z(n14686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6144_3_lut.init = 16'hcaca;
    LUT4 i6113_3_lut (.A(n14653), .B(n14654), .C(r_addr[4]), .Z(n14655)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6113_3_lut.init = 16'hcaca;
    LUT4 i6082_3_lut (.A(n14622), .B(n14623), .C(r_addr[4]), .Z(n14624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6082_3_lut.init = 16'hcaca;
    LUT4 i6051_3_lut (.A(n14591), .B(n14592), .C(r_addr[4]), .Z(n14593)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6051_3_lut.init = 16'hcaca;
    LUT4 i6020_3_lut (.A(n14560), .B(n14561), .C(r_addr[4]), .Z(n14562)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6020_3_lut.init = 16'hcaca;
    LUT4 i5989_3_lut (.A(n14529), .B(n14530), .C(r_addr[4]), .Z(n14531)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5989_3_lut.init = 16'hcaca;
    LUT4 i5124_3_lut (.A(n13664), .B(n13665), .C(r_addr[4]), .Z(n13666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5124_3_lut.init = 16'hcaca;
    LUT4 i5093_3_lut (.A(n13633), .B(n13634), .C(r_addr[4]), .Z(n13635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5093_3_lut.init = 16'hcaca;
    LUT4 i5062_3_lut (.A(n13602), .B(n13603), .C(r_addr[4]), .Z(n13604)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5062_3_lut.init = 16'hcaca;
    LUT4 i5031_3_lut (.A(n13571), .B(n13572), .C(r_addr[4]), .Z(n13573)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5031_3_lut.init = 16'hcaca;
    LUT4 i5000_3_lut (.A(n13540), .B(n13541), .C(r_addr[4]), .Z(n13542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5000_3_lut.init = 16'hcaca;
    LUT4 i4969_3_lut (.A(n13509), .B(n13510), .C(r_addr[4]), .Z(n13511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4969_3_lut.init = 16'hcaca;
    LUT4 i4869_3_lut (.A(n13409), .B(n13410), .C(r_addr[4]), .Z(n13411)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4869_3_lut.init = 16'hcaca;
    LUT4 i4838_3_lut (.A(n13378), .B(n13379), .C(r_addr[4]), .Z(n13380)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4838_3_lut.init = 16'hcaca;
    LUT4 i4807_3_lut (.A(n13347), .B(n13348), .C(r_addr[4]), .Z(n13349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4807_3_lut.init = 16'hcaca;
    LUT4 i4776_3_lut (.A(n13316), .B(n13317), .C(r_addr[4]), .Z(n13318)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4776_3_lut.init = 16'hcaca;
    LUT4 i4745_3_lut (.A(n13285), .B(n13286), .C(r_addr[4]), .Z(n13287)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4745_3_lut.init = 16'hcaca;
    LUT4 i4714_3_lut (.A(n13254), .B(n13255), .C(r_addr[4]), .Z(n13256)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4714_3_lut.init = 16'hcaca;
    LUT4 i5634_3_lut (.A(n14174), .B(n14175), .C(r_addr[4]), .Z(n14176)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5634_3_lut.init = 16'hcaca;
    LUT4 i5603_3_lut (.A(n14143), .B(n14144), .C(r_addr[4]), .Z(n14145)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5603_3_lut.init = 16'hcaca;
    LUT4 i5572_3_lut (.A(n14112), .B(n14113), .C(r_addr[4]), .Z(n14114)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5572_3_lut.init = 16'hcaca;
    LUT4 i5541_3_lut (.A(n14081), .B(n14082), .C(r_addr[4]), .Z(n14083)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5541_3_lut.init = 16'hcaca;
    LUT4 i5510_3_lut (.A(n14050), .B(n14051), .C(r_addr[4]), .Z(n14052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5510_3_lut.init = 16'hcaca;
    LUT4 i5479_3_lut (.A(n14019), .B(n14020), .C(r_addr[4]), .Z(n14021)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5479_3_lut.init = 16'hcaca;
    LUT4 i6399_3_lut (.A(n14939), .B(n14940), .C(r_addr[4]), .Z(n14941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6399_3_lut.init = 16'hcaca;
    LUT4 i6368_3_lut (.A(n14908), .B(n14909), .C(r_addr[4]), .Z(n14910)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6368_3_lut.init = 16'hcaca;
    LUT4 i4614_3_lut (.A(n13154), .B(n13155), .C(r_addr[4]), .Z(n13156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4614_3_lut.init = 16'hcaca;
    LUT4 i4583_3_lut (.A(n13123), .B(n13124), .C(r_addr[4]), .Z(n13125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4583_3_lut.init = 16'hcaca;
    LUT4 i4552_3_lut (.A(n13092), .B(n13093), .C(r_addr[4]), .Z(n13094)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4552_3_lut.init = 16'hcaca;
    LUT4 i4521_3_lut (.A(n13061), .B(n13062), .C(r_addr[4]), .Z(n13063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4521_3_lut.init = 16'hcaca;
    LUT4 i4490_3_lut (.A(n13030), .B(n13031), .C(r_addr[4]), .Z(n13032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4490_3_lut.init = 16'hcaca;
    LUT4 i4459_3_lut (.A(n12999), .B(n13000), .C(r_addr[4]), .Z(n13001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4459_3_lut.init = 16'hcaca;
    LUT4 i6337_3_lut (.A(n14877), .B(n14878), .C(r_addr[4]), .Z(n14879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6337_3_lut.init = 16'hcaca;
    LUT4 i6306_3_lut (.A(n14846), .B(n14847), .C(r_addr[4]), .Z(n14848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6306_3_lut.init = 16'hcaca;
    LUT4 i4428_3_lut (.A(n12968), .B(n12969), .C(r_addr[4]), .Z(n12970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4428_3_lut.init = 16'hcaca;
    LUT4 i4397_3_lut (.A(n12937), .B(n12938), .C(r_addr[4]), .Z(n12939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4397_3_lut.init = 16'hcaca;
    LUT4 i4683_3_lut (.A(n13223), .B(n13224), .C(r_addr[4]), .Z(n13225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4683_3_lut.init = 16'hcaca;
    LUT4 i4652_3_lut (.A(n13192), .B(n13193), .C(r_addr[4]), .Z(n13194)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4652_3_lut.init = 16'hcaca;
    LUT4 i4938_3_lut (.A(n13478), .B(n13479), .C(r_addr[4]), .Z(n13480)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4938_3_lut.init = 16'hcaca;
    LUT4 i4907_3_lut (.A(n13447), .B(n13448), .C(r_addr[4]), .Z(n13449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i4907_3_lut.init = 16'hcaca;
    LUT4 i5193_3_lut (.A(n13733), .B(n13734), .C(r_addr[4]), .Z(n13735)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5193_3_lut.init = 16'hcaca;
    LUT4 i5162_3_lut (.A(n13702), .B(n13703), .C(r_addr[4]), .Z(n13704)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5162_3_lut.init = 16'hcaca;
    LUT4 i5448_3_lut (.A(n13988), .B(n13989), .C(r_addr[4]), .Z(n13990)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5448_3_lut.init = 16'hcaca;
    LUT4 i5417_3_lut (.A(n13957), .B(n13958), .C(r_addr[4]), .Z(n13959)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5417_3_lut.init = 16'hcaca;
    LUT4 i5703_3_lut (.A(n14243), .B(n14244), .C(r_addr[4]), .Z(n14245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5703_3_lut.init = 16'hcaca;
    LUT4 i5672_3_lut (.A(n14212), .B(n14213), .C(r_addr[4]), .Z(n14214)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5672_3_lut.init = 16'hcaca;
    LUT4 i5958_3_lut (.A(n14498), .B(n14499), .C(r_addr[4]), .Z(n14500)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5958_3_lut.init = 16'hcaca;
    LUT4 i5927_3_lut (.A(n14467), .B(n14468), .C(r_addr[4]), .Z(n14469)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5927_3_lut.init = 16'hcaca;
    LUT4 i6213_3_lut (.A(n14753), .B(n14754), .C(r_addr[4]), .Z(n14755)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6213_3_lut.init = 16'hcaca;
    LUT4 i6182_3_lut (.A(n14722), .B(n14723), .C(r_addr[4]), .Z(n14724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6182_3_lut.init = 16'hcaca;
    LUT4 i6275_3_lut (.A(n14815), .B(n14816), .C(r_addr[4]), .Z(n14817)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6275_3_lut.init = 16'hcaca;
    LUT4 i6244_3_lut (.A(n14784), .B(n14785), .C(r_addr[4]), .Z(n14786)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6244_3_lut.init = 16'hcaca;
    LUT4 i5379_3_lut (.A(n13919), .B(n13920), .C(r_addr[4]), .Z(n13921)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5379_3_lut.init = 16'hcaca;
    LUT4 i5348_3_lut (.A(n13888), .B(n13889), .C(r_addr[4]), .Z(n13890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5348_3_lut.init = 16'hcaca;
    LUT4 i5317_3_lut (.A(n13857), .B(n13858), .C(r_addr[4]), .Z(n13859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5317_3_lut.init = 16'hcaca;
    LUT4 i5286_3_lut (.A(n13826), .B(n13827), .C(r_addr[4]), .Z(n13828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5286_3_lut.init = 16'hcaca;
    LUT4 i5255_3_lut (.A(n13795), .B(n13796), .C(r_addr[4]), .Z(n13797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5255_3_lut.init = 16'hcaca;
    LUT4 i5224_3_lut (.A(n13764), .B(n13765), .C(r_addr[4]), .Z(n13766)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5224_3_lut.init = 16'hcaca;
    LUT4 i5889_3_lut (.A(n14429), .B(n14430), .C(r_addr[4]), .Z(n14431)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5889_3_lut.init = 16'hcaca;
    LUT4 i5858_3_lut (.A(n14398), .B(n14399), .C(r_addr[4]), .Z(n14400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5858_3_lut.init = 16'hcaca;
    LUT4 i5827_3_lut (.A(n14367), .B(n14368), .C(r_addr[4]), .Z(n14369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5827_3_lut.init = 16'hcaca;
    LUT4 i5796_3_lut (.A(n14336), .B(n14337), .C(r_addr[4]), .Z(n14338)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5796_3_lut.init = 16'hcaca;
    LUT4 i5765_3_lut (.A(n14305), .B(n14306), .C(r_addr[4]), .Z(n14307)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5765_3_lut.init = 16'hcaca;
    LUT4 i5734_3_lut (.A(n14274), .B(n14275), .C(r_addr[4]), .Z(n14276)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5734_3_lut.init = 16'hcaca;
    LUT4 i787_2_lut (.A(rd_en_c), .B(clk_c_enable_1007), .Z(clk_c_enable_2057)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(33[12] 36[12])
    defparam i787_2_lut.init = 16'h2222;
    LUT4 mux_220_i2_3_lut_4_lut (.A(n15014), .B(n14994), .C(\array[39] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2369[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_220_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_220_i3_3_lut_4_lut (.A(n15014), .B(n14994), .C(\array[39] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2369[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_220_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_220_i4_3_lut_4_lut (.A(n15014), .B(n14994), .C(\array[39] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2369[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_220_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_220_i5_3_lut_4_lut (.A(n15014), .B(n14994), .C(\array[39] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2369[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_220_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_220_i6_3_lut_4_lut (.A(n15014), .B(n14994), .C(\array[39] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2369[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_220_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_220_i7_3_lut_4_lut (.A(n15014), .B(n14994), .C(\array[39] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2369[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_220_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_220_i8_3_lut_4_lut (.A(n15014), .B(n14994), .C(\array[39] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2369[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_220_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_259_i1_3_lut_4_lut (.A(n15007), .B(n14992), .C(\array[0] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2057[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_259_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_259_i2_3_lut_4_lut (.A(n15007), .B(n14992), .C(\array[0] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2057[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_259_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_259_i3_3_lut_4_lut (.A(n15007), .B(n14992), .C(\array[0] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2057[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_259_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_259_i4_3_lut_4_lut (.A(n15007), .B(n14992), .C(\array[0] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2057[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_259_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_259_i5_3_lut_4_lut (.A(n15007), .B(n14992), .C(\array[0] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2057[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_259_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_259_i6_3_lut_4_lut (.A(n15007), .B(n14992), .C(\array[0] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2057[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_259_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_259_i7_3_lut_4_lut (.A(n15007), .B(n14992), .C(\array[0] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2057[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_259_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_259_i8_3_lut_4_lut (.A(n15007), .B(n14992), .C(\array[0] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2057[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_259_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_258_i1_3_lut_4_lut (.A(n15008), .B(n14992), .C(\array[1] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2065[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_258_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_258_i2_3_lut_4_lut (.A(n15008), .B(n14992), .C(\array[1] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2065[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_258_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_258_i3_3_lut_4_lut (.A(n15008), .B(n14992), .C(\array[1] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2065[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_258_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_258_i4_3_lut_4_lut (.A(n15008), .B(n14992), .C(\array[1] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2065[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_258_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_258_i5_3_lut_4_lut (.A(n15008), .B(n14992), .C(\array[1] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2065[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_258_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_258_i6_3_lut_4_lut (.A(n15008), .B(n14992), .C(\array[1] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2065[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_258_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_258_i7_3_lut_4_lut (.A(n15008), .B(n14992), .C(\array[1] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2065[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_258_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_258_i8_3_lut_4_lut (.A(n15008), .B(n14992), .C(\array[1] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2065[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_258_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_257_i1_3_lut_4_lut (.A(n15009), .B(n14992), .C(\array[2] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2073[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_257_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_257_i2_3_lut_4_lut (.A(n15009), .B(n14992), .C(\array[2] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2073[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_257_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_257_i3_3_lut_4_lut (.A(n15009), .B(n14992), .C(\array[2] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2073[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_257_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5333_3_lut (.A(\array[222] [4]), .B(\array[223] [4]), .C(r_addr[0]), 
         .Z(n13875)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5333_3_lut.init = 16'hcaca;
    LUT4 i5332_3_lut (.A(\array[220] [4]), .B(\array[221] [4]), .C(r_addr[0]), 
         .Z(n13874)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5332_3_lut.init = 16'hcaca;
    LUT4 mux_257_i4_3_lut_4_lut (.A(n15009), .B(n14992), .C(\array[2] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2073[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_257_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_257_i5_3_lut_4_lut (.A(n15009), .B(n14992), .C(\array[2] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2073[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_257_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5874_3_lut (.A(\array[254] [6]), .B(\array[255] [6]), .C(r_addr[0]), 
         .Z(n14416)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5874_3_lut.init = 16'hcaca;
    LUT4 i5873_3_lut (.A(\array[252] [6]), .B(\array[253] [6]), .C(r_addr[0]), 
         .Z(n14415)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5873_3_lut.init = 16'hcaca;
    LUT4 i5331_3_lut (.A(\array[218] [4]), .B(\array[219] [4]), .C(r_addr[0]), 
         .Z(n13873)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5331_3_lut.init = 16'hcaca;
    LUT4 mux_257_i6_3_lut_4_lut (.A(n15009), .B(n14992), .C(\array[2] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2073[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_257_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_257_i7_3_lut_4_lut (.A(n15009), .B(n14992), .C(\array[2] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2073[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_257_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_257_i8_3_lut_4_lut (.A(n15009), .B(n14992), .C(\array[2] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2073[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_257_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_256_i1_3_lut_4_lut (.A(n15010), .B(n14992), .C(\array[3] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2081[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_256_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_256_i2_3_lut_4_lut (.A(n15010), .B(n14992), .C(\array[3] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2081[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_256_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_256_i3_3_lut_4_lut (.A(n15010), .B(n14992), .C(\array[3] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2081[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_256_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_256_i4_3_lut_4_lut (.A(n15010), .B(n14992), .C(\array[3] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2081[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_256_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_256_i5_3_lut_4_lut (.A(n15010), .B(n14992), .C(\array[3] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2081[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_256_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_256_i6_3_lut_4_lut (.A(n15010), .B(n14992), .C(\array[3] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2081[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_256_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_256_i7_3_lut_4_lut (.A(n15010), .B(n14992), .C(\array[3] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2081[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_256_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_256_i8_3_lut_4_lut (.A(n15010), .B(n14992), .C(\array[3] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2081[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_256_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5330_3_lut (.A(\array[216] [4]), .B(\array[217] [4]), .C(r_addr[0]), 
         .Z(n13872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i5330_3_lut.init = 16'hcaca;
    LUT4 mux_255_i1_3_lut_4_lut (.A(n15011), .B(n14992), .C(\array[4] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2089[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_255_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_255_i2_3_lut_4_lut (.A(n15011), .B(n14992), .C(\array[4] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2089[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_255_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_252_i3_3_lut_4_lut (.A(n15014), .B(n14992), .C(\array[7] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2113[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_252_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_252_i4_3_lut_4_lut (.A(n15014), .B(n14992), .C(\array[7] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2113[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_252_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_252_i5_3_lut_4_lut (.A(n15014), .B(n14992), .C(\array[7] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2113[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_252_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_252_i6_3_lut_4_lut (.A(n15014), .B(n14992), .C(\array[7] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2113[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_252_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_252_i7_3_lut_4_lut (.A(n15014), .B(n14992), .C(\array[7] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2113[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_252_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_252_i8_3_lut_4_lut (.A(n15014), .B(n14992), .C(\array[7] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2113[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_252_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_251_i1_3_lut_4_lut (.A(n15015), .B(n14992), .C(\array[8] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2121[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_251_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_251_i2_3_lut_4_lut (.A(n15015), .B(n14992), .C(\array[8] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2121[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_251_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_251_i3_3_lut_4_lut (.A(n15015), .B(n14992), .C(\array[8] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2121[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_251_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_251_i4_3_lut_4_lut (.A(n15015), .B(n14992), .C(\array[8] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2121[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_251_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_251_i5_3_lut_4_lut (.A(n15015), .B(n14992), .C(\array[8] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2121[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_251_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_251_i6_3_lut_4_lut (.A(n15015), .B(n14992), .C(\array[8] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2121[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_251_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_251_i7_3_lut_4_lut (.A(n15015), .B(n14992), .C(\array[8] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2121[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_251_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_251_i8_3_lut_4_lut (.A(n15015), .B(n14992), .C(\array[8] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2121[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_251_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_250_i1_3_lut_4_lut (.A(n15016), .B(n14992), .C(\array[9] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2129[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_250_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_250_i2_3_lut_4_lut (.A(n15016), .B(n14992), .C(\array[9] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2129[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_250_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_250_i3_3_lut_4_lut (.A(n15016), .B(n14992), .C(\array[9] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2129[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_250_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_250_i4_3_lut_4_lut (.A(n15016), .B(n14992), .C(\array[9] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2129[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_250_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_250_i5_3_lut_4_lut (.A(n15016), .B(n14992), .C(\array[9] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2129[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_250_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_250_i6_3_lut_4_lut (.A(n15016), .B(n14992), .C(\array[9] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2129[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_250_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_250_i7_3_lut_4_lut (.A(n15016), .B(n14992), .C(\array[9] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2129[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_250_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_250_i8_3_lut_4_lut (.A(n15016), .B(n14992), .C(\array[9] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2129[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_250_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_249_i1_3_lut_4_lut (.A(n15017), .B(n14992), .C(\array[10] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2137[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_249_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_249_i2_3_lut_4_lut (.A(n15017), .B(n14992), .C(\array[10] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2137[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_249_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_249_i3_3_lut_4_lut (.A(n15017), .B(n14992), .C(\array[10] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2137[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_249_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_249_i4_3_lut_4_lut (.A(n15017), .B(n14992), .C(\array[10] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2137[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_249_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_249_i5_3_lut_4_lut (.A(n15017), .B(n14992), .C(\array[10] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2137[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_249_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_249_i6_3_lut_4_lut (.A(n15017), .B(n14992), .C(\array[10] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2137[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_249_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_249_i7_3_lut_4_lut (.A(n15017), .B(n14992), .C(\array[10] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2137[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_249_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_249_i8_3_lut_4_lut (.A(n15017), .B(n14992), .C(\array[10] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2137[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_249_i8_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX r_addr_i0_i1 (.D(addr_c_1), .SP(clk_c_enable_2057), .CK(clk_c), 
            .Q(r_addr[1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam r_addr_i0_i1.GSR = "ENABLED";
    GSR GSR_INST (.GSR(VCC_net));
    LUT4 mux_248_i1_3_lut_4_lut (.A(n15018), .B(n14992), .C(\array[11] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2145[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_248_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_248_i2_3_lut_4_lut (.A(n15018), .B(n14992), .C(\array[11] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2145[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_248_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_248_i3_3_lut_4_lut (.A(n15018), .B(n14992), .C(\array[11] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2145[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_248_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_248_i4_3_lut_4_lut (.A(n15018), .B(n14992), .C(\array[11] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2145[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_248_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_248_i5_3_lut_4_lut (.A(n15018), .B(n14992), .C(\array[11] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2145[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_248_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_248_i6_3_lut_4_lut (.A(n15018), .B(n14992), .C(\array[11] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2145[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_248_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_248_i7_3_lut_4_lut (.A(n15018), .B(n14992), .C(\array[11] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2145[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_248_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_248_i8_3_lut_4_lut (.A(n15018), .B(n14992), .C(\array[11] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2145[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_248_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_247_i1_3_lut_4_lut (.A(n15019), .B(n14992), .C(\array[12] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2153[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_247_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_247_i2_3_lut_4_lut (.A(n15019), .B(n14992), .C(\array[12] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2153[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_247_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_247_i3_3_lut_4_lut (.A(n15019), .B(n14992), .C(\array[12] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2153[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_247_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_247_i4_3_lut_4_lut (.A(n15019), .B(n14992), .C(\array[12] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2153[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_247_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_247_i5_3_lut_4_lut (.A(n15019), .B(n14992), .C(\array[12] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2153[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_247_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_247_i6_3_lut_4_lut (.A(n15019), .B(n14992), .C(\array[12] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2153[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_247_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_247_i7_3_lut_4_lut (.A(n15019), .B(n14992), .C(\array[12] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2153[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_247_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_247_i8_3_lut_4_lut (.A(n15019), .B(n14992), .C(\array[12] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2153[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_247_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_246_i1_3_lut_4_lut (.A(n15020), .B(n14992), .C(\array[13] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2161[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_246_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_246_i2_3_lut_4_lut (.A(n15020), .B(n14992), .C(\array[13] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2161[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_246_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_246_i3_3_lut_4_lut (.A(n15020), .B(n14992), .C(\array[13] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2161[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_246_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_246_i4_3_lut_4_lut (.A(n15020), .B(n14992), .C(\array[13] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2161[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_246_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_246_i5_3_lut_4_lut (.A(n15020), .B(n14992), .C(\array[13] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2161[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_246_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_246_i6_3_lut_4_lut (.A(n15020), .B(n14992), .C(\array[13] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2161[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_246_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_246_i7_3_lut_4_lut (.A(n15020), .B(n14992), .C(\array[13] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2161[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_246_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_246_i8_3_lut_4_lut (.A(n15020), .B(n14992), .C(\array[13] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2161[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_246_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_245_i1_3_lut_4_lut (.A(n15021), .B(n14992), .C(\array[14] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2169[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_245_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_245_i2_3_lut_4_lut (.A(n15021), .B(n14992), .C(\array[14] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2169[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_245_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_245_i3_3_lut_4_lut (.A(n15021), .B(n14992), .C(\array[14] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2169[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_245_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_245_i4_3_lut_4_lut (.A(n15021), .B(n14992), .C(\array[14] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2169[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_245_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_245_i5_3_lut_4_lut (.A(n15021), .B(n14992), .C(\array[14] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2169[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_245_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_245_i6_3_lut_4_lut (.A(n15021), .B(n14992), .C(\array[14] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2169[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_245_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_245_i7_3_lut_4_lut (.A(n15021), .B(n14992), .C(\array[14] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2169[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_245_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_245_i8_3_lut_4_lut (.A(n15021), .B(n14992), .C(\array[14] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2169[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_245_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_244_i1_3_lut_4_lut (.A(n15023), .B(n14992), .C(\array[15] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2177[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_244_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_244_i2_3_lut_4_lut (.A(n15023), .B(n14992), .C(\array[15] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2177[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_244_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_244_i3_3_lut_4_lut (.A(n15023), .B(n14992), .C(\array[15] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2177[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_244_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_244_i4_3_lut_4_lut (.A(n15023), .B(n14992), .C(\array[15] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2177[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_244_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_244_i5_3_lut_4_lut (.A(n15023), .B(n14992), .C(\array[15] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2177[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_244_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_244_i6_3_lut_4_lut (.A(n15023), .B(n14992), .C(\array[15] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2177[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_244_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_244_i7_3_lut_4_lut (.A(n15023), .B(n14992), .C(\array[15] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2177[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_244_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_244_i8_3_lut_4_lut (.A(n15023), .B(n14992), .C(\array[15] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2177[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_244_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_243_i1_3_lut_4_lut (.A(n15007), .B(n14993), .C(\array[16] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2185[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_243_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_243_i2_3_lut_4_lut (.A(n15007), .B(n14993), .C(\array[16] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2185[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_243_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_243_i3_3_lut_4_lut (.A(n15007), .B(n14993), .C(\array[16] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2185[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_243_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_243_i4_3_lut_4_lut (.A(n15007), .B(n14993), .C(\array[16] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2185[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_243_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_243_i5_3_lut_4_lut (.A(n15007), .B(n14993), .C(\array[16] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2185[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_243_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_243_i6_3_lut_4_lut (.A(n15007), .B(n14993), .C(\array[16] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2185[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_243_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_243_i7_3_lut_4_lut (.A(n15007), .B(n14993), .C(\array[16] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2185[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_243_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_243_i8_3_lut_4_lut (.A(n15007), .B(n14993), .C(\array[16] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2185[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_243_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_242_i1_3_lut_4_lut (.A(n15008), .B(n14993), .C(\array[17] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2193[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_242_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_242_i2_3_lut_4_lut (.A(n15008), .B(n14993), .C(\array[17] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2193[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_242_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_242_i3_3_lut_4_lut (.A(n15008), .B(n14993), .C(\array[17] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2193[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_242_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_242_i4_3_lut_4_lut (.A(n15008), .B(n14993), .C(\array[17] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2193[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_242_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_242_i5_3_lut_4_lut (.A(n15008), .B(n14993), .C(\array[17] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2193[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_242_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_242_i6_3_lut_4_lut (.A(n15008), .B(n14993), .C(\array[17] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2193[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_242_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_242_i7_3_lut_4_lut (.A(n15008), .B(n14993), .C(\array[17] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2193[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_242_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_242_i8_3_lut_4_lut (.A(n15008), .B(n14993), .C(\array[17] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2193[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_242_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_241_i1_3_lut_4_lut (.A(n15009), .B(n14993), .C(\array[18] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2201[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_241_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_241_i2_3_lut_4_lut (.A(n15009), .B(n14993), .C(\array[18] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2201[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_241_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_241_i3_3_lut_4_lut (.A(n15009), .B(n14993), .C(\array[18] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2201[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_241_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_241_i4_3_lut_4_lut (.A(n15009), .B(n14993), .C(\array[18] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2201[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_241_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_241_i5_3_lut_4_lut (.A(n15009), .B(n14993), .C(\array[18] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2201[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_241_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_241_i6_3_lut_4_lut (.A(n15009), .B(n14993), .C(\array[18] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2201[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_241_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_241_i7_3_lut_4_lut (.A(n15009), .B(n14993), .C(\array[18] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2201[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_241_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_241_i8_3_lut_4_lut (.A(n15009), .B(n14993), .C(\array[18] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2201[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_241_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_240_i1_3_lut_4_lut (.A(n15010), .B(n14993), .C(\array[19] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2209[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_240_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_240_i2_3_lut_4_lut (.A(n15010), .B(n14993), .C(\array[19] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2209[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_240_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_240_i3_3_lut_4_lut (.A(n15010), .B(n14993), .C(\array[19] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2209[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_240_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_240_i4_3_lut_4_lut (.A(n15010), .B(n14993), .C(\array[19] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2209[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_240_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_240_i5_3_lut_4_lut (.A(n15010), .B(n14993), .C(\array[19] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2209[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_240_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_240_i6_3_lut_4_lut (.A(n15010), .B(n14993), .C(\array[19] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2209[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_240_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_240_i7_3_lut_4_lut (.A(n15010), .B(n14993), .C(\array[19] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2209[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_240_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_240_i8_3_lut_4_lut (.A(n15010), .B(n14993), .C(\array[19] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2209[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_240_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_239_i1_3_lut_4_lut (.A(n15011), .B(n14993), .C(\array[20] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2217[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_239_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_239_i2_3_lut_4_lut (.A(n15011), .B(n14993), .C(\array[20] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2217[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_239_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_239_i3_3_lut_4_lut (.A(n15011), .B(n14993), .C(\array[20] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2217[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_239_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_239_i4_3_lut_4_lut (.A(n15011), .B(n14993), .C(\array[20] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2217[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_239_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_239_i5_3_lut_4_lut (.A(n15011), .B(n14993), .C(\array[20] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2217[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_239_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_239_i6_3_lut_4_lut (.A(n15011), .B(n14993), .C(\array[20] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2217[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_239_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_239_i7_3_lut_4_lut (.A(n15011), .B(n14993), .C(\array[20] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2217[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_239_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_239_i8_3_lut_4_lut (.A(n15011), .B(n14993), .C(\array[20] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2217[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_239_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_238_i1_3_lut_4_lut (.A(n15012), .B(n14993), .C(\array[21] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2225[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_238_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_238_i2_3_lut_4_lut (.A(n15012), .B(n14993), .C(\array[21] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2225[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_238_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_238_i3_3_lut_4_lut (.A(n15012), .B(n14993), .C(\array[21] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2225[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_238_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_238_i4_3_lut_4_lut (.A(n15012), .B(n14993), .C(\array[21] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2225[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_238_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_238_i5_3_lut_4_lut (.A(n15012), .B(n14993), .C(\array[21] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2225[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_238_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_238_i6_3_lut_4_lut (.A(n15012), .B(n14993), .C(\array[21] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2225[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_238_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_238_i7_3_lut_4_lut (.A(n15012), .B(n14993), .C(\array[21] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2225[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_238_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_238_i8_3_lut_4_lut (.A(n15012), .B(n14993), .C(\array[21] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2225[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_238_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_237_i1_3_lut_4_lut (.A(n15013), .B(n14993), .C(\array[22] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2233[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_237_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_237_i2_3_lut_4_lut (.A(n15013), .B(n14993), .C(\array[22] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2233[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_237_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_237_i3_3_lut_4_lut (.A(n15013), .B(n14993), .C(\array[22] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2233[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_237_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_237_i4_3_lut_4_lut (.A(n15013), .B(n14993), .C(\array[22] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2233[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_237_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_237_i5_3_lut_4_lut (.A(n15013), .B(n14993), .C(\array[22] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2233[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_237_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_237_i6_3_lut_4_lut (.A(n15013), .B(n14993), .C(\array[22] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2233[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_237_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_237_i7_3_lut_4_lut (.A(n15013), .B(n14993), .C(\array[22] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2233[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_237_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_237_i8_3_lut_4_lut (.A(n15013), .B(n14993), .C(\array[22] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2233[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_237_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_236_i1_3_lut_4_lut (.A(n15014), .B(n14993), .C(\array[23] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2241[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_236_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_236_i2_3_lut_4_lut (.A(n15014), .B(n14993), .C(\array[23] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2241[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_236_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_236_i3_3_lut_4_lut (.A(n15014), .B(n14993), .C(\array[23] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2241[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_236_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_236_i4_3_lut_4_lut (.A(n15014), .B(n14993), .C(\array[23] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2241[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_236_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_236_i5_3_lut_4_lut (.A(n15014), .B(n14993), .C(\array[23] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2241[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_236_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_236_i6_3_lut_4_lut (.A(n15014), .B(n14993), .C(\array[23] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2241[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_236_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_236_i7_3_lut_4_lut (.A(n15014), .B(n14993), .C(\array[23] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2241[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_236_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_236_i8_3_lut_4_lut (.A(n15014), .B(n14993), .C(\array[23] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2241[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_236_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_235_i1_3_lut_4_lut (.A(n15015), .B(n14993), .C(\array[24] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2249[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_235_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_235_i2_3_lut_4_lut (.A(n15015), .B(n14993), .C(\array[24] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2249[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_235_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_235_i3_3_lut_4_lut (.A(n15015), .B(n14993), .C(\array[24] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2249[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_235_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_235_i4_3_lut_4_lut (.A(n15015), .B(n14993), .C(\array[24] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2249[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_235_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_235_i5_3_lut_4_lut (.A(n15015), .B(n14993), .C(\array[24] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2249[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_235_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_235_i6_3_lut_4_lut (.A(n15015), .B(n14993), .C(\array[24] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2249[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_235_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_235_i7_3_lut_4_lut (.A(n15015), .B(n14993), .C(\array[24] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2249[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_235_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_235_i8_3_lut_4_lut (.A(n15015), .B(n14993), .C(\array[24] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2249[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_235_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_234_i1_3_lut_4_lut (.A(n15016), .B(n14993), .C(\array[25] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2257[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_234_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_234_i2_3_lut_4_lut (.A(n15016), .B(n14993), .C(\array[25] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2257[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_234_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_234_i3_3_lut_4_lut (.A(n15016), .B(n14993), .C(\array[25] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2257[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_234_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_234_i4_3_lut_4_lut (.A(n15016), .B(n14993), .C(\array[25] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2257[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_234_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_234_i5_3_lut_4_lut (.A(n15016), .B(n14993), .C(\array[25] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2257[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_234_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_234_i6_3_lut_4_lut (.A(n15016), .B(n14993), .C(\array[25] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2257[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_234_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_234_i7_3_lut_4_lut (.A(n15016), .B(n14993), .C(\array[25] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2257[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_234_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_234_i8_3_lut_4_lut (.A(n15016), .B(n14993), .C(\array[25] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2257[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_234_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_233_i1_3_lut_4_lut (.A(n15017), .B(n14993), .C(\array[26] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2265[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_233_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_233_i2_3_lut_4_lut (.A(n15017), .B(n14993), .C(\array[26] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2265[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_233_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_233_i3_3_lut_4_lut (.A(n15017), .B(n14993), .C(\array[26] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2265[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_233_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_233_i4_3_lut_4_lut (.A(n15017), .B(n14993), .C(\array[26] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2265[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_233_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_233_i5_3_lut_4_lut (.A(n15017), .B(n14993), .C(\array[26] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2265[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_233_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_233_i6_3_lut_4_lut (.A(n15017), .B(n14993), .C(\array[26] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2265[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_233_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_233_i7_3_lut_4_lut (.A(n15017), .B(n14993), .C(\array[26] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2265[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_233_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_233_i8_3_lut_4_lut (.A(n15017), .B(n14993), .C(\array[26] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2265[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_233_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_232_i1_3_lut_4_lut (.A(n15018), .B(n14993), .C(\array[27] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2273[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_232_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_255_i3_3_lut_4_lut (.A(n15011), .B(n14992), .C(\array[4] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2089[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_255_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_232_i2_3_lut_4_lut (.A(n15018), .B(n14993), .C(\array[27] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2273[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_232_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_232_i3_3_lut_4_lut (.A(n15018), .B(n14993), .C(\array[27] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2273[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_232_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_232_i4_3_lut_4_lut (.A(n15018), .B(n14993), .C(\array[27] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2273[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_232_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_232_i5_3_lut_4_lut (.A(n15018), .B(n14993), .C(\array[27] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2273[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_232_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_232_i6_3_lut_4_lut (.A(n15018), .B(n14993), .C(\array[27] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2273[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_232_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_232_i7_3_lut_4_lut (.A(n15018), .B(n14993), .C(\array[27] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2273[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_232_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_232_i8_3_lut_4_lut (.A(n15018), .B(n14993), .C(\array[27] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2273[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_232_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_231_i1_3_lut_4_lut (.A(n15019), .B(n14993), .C(\array[28] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2281[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_231_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_231_i2_3_lut_4_lut (.A(n15019), .B(n14993), .C(\array[28] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2281[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_231_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_231_i3_3_lut_4_lut (.A(n15019), .B(n14993), .C(\array[28] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2281[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_231_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_231_i4_3_lut_4_lut (.A(n15019), .B(n14993), .C(\array[28] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2281[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_231_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_231_i5_3_lut_4_lut (.A(n15019), .B(n14993), .C(\array[28] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2281[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_231_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_231_i6_3_lut_4_lut (.A(n15019), .B(n14993), .C(\array[28] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2281[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_231_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_231_i7_3_lut_4_lut (.A(n15019), .B(n14993), .C(\array[28] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2281[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_231_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_231_i8_3_lut_4_lut (.A(n15019), .B(n14993), .C(\array[28] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2281[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_231_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_230_i1_3_lut_4_lut (.A(n15020), .B(n14993), .C(\array[29] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2289[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_230_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_230_i2_3_lut_4_lut (.A(n15020), .B(n14993), .C(\array[29] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2289[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_230_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_230_i3_3_lut_4_lut (.A(n15020), .B(n14993), .C(\array[29] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2289[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_230_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_230_i4_3_lut_4_lut (.A(n15020), .B(n14993), .C(\array[29] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2289[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_230_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_230_i5_3_lut_4_lut (.A(n15020), .B(n14993), .C(\array[29] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2289[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_230_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_230_i6_3_lut_4_lut (.A(n15020), .B(n14993), .C(\array[29] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2289[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_230_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_230_i7_3_lut_4_lut (.A(n15020), .B(n14993), .C(\array[29] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2289[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_230_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_230_i8_3_lut_4_lut (.A(n15020), .B(n14993), .C(\array[29] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2289[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_230_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_229_i1_3_lut_4_lut (.A(n15021), .B(n14993), .C(\array[30] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2297[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_229_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_229_i2_3_lut_4_lut (.A(n15021), .B(n14993), .C(\array[30] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2297[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_229_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_229_i3_3_lut_4_lut (.A(n15021), .B(n14993), .C(\array[30] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2297[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_229_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_229_i4_3_lut_4_lut (.A(n15021), .B(n14993), .C(\array[30] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2297[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_229_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_229_i5_3_lut_4_lut (.A(n15021), .B(n14993), .C(\array[30] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2297[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_229_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_229_i6_3_lut_4_lut (.A(n15021), .B(n14993), .C(\array[30] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2297[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_229_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_229_i7_3_lut_4_lut (.A(n15021), .B(n14993), .C(\array[30] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2297[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_229_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_229_i8_3_lut_4_lut (.A(n15021), .B(n14993), .C(\array[30] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2297[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_229_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_228_i1_3_lut_4_lut (.A(n15023), .B(n14993), .C(\array[31] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2305[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_228_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_228_i2_3_lut_4_lut (.A(n15023), .B(n14993), .C(\array[31] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2305[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_228_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_228_i3_3_lut_4_lut (.A(n15023), .B(n14993), .C(\array[31] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2305[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_228_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_228_i4_3_lut_4_lut (.A(n15023), .B(n14993), .C(\array[31] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2305[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_228_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_228_i5_3_lut_4_lut (.A(n15023), .B(n14993), .C(\array[31] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2305[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_228_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_228_i6_3_lut_4_lut (.A(n15023), .B(n14993), .C(\array[31] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2305[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_228_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_228_i7_3_lut_4_lut (.A(n15023), .B(n14993), .C(\array[31] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2305[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_228_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_228_i8_3_lut_4_lut (.A(n15023), .B(n14993), .C(\array[31] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2305[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_228_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_227_i1_3_lut_4_lut (.A(n15007), .B(n14994), .C(\array[32] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2313[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_227_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_227_i2_3_lut_4_lut (.A(n15007), .B(n14994), .C(\array[32] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2313[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_227_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_227_i3_3_lut_4_lut (.A(n15007), .B(n14994), .C(\array[32] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2313[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_227_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_227_i4_3_lut_4_lut (.A(n15007), .B(n14994), .C(\array[32] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2313[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_227_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_227_i5_3_lut_4_lut (.A(n15007), .B(n14994), .C(\array[32] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2313[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_227_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_227_i6_3_lut_4_lut (.A(n15007), .B(n14994), .C(\array[32] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2313[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_227_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_227_i7_3_lut_4_lut (.A(n15007), .B(n14994), .C(\array[32] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2313[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_227_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_227_i8_3_lut_4_lut (.A(n15007), .B(n14994), .C(\array[32] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2313[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_227_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_226_i1_3_lut_4_lut (.A(n15008), .B(n14994), .C(\array[33] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2321[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_226_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_226_i2_3_lut_4_lut (.A(n15008), .B(n14994), .C(\array[33] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2321[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_226_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_226_i3_3_lut_4_lut (.A(n15008), .B(n14994), .C(\array[33] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2321[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_226_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_226_i4_3_lut_4_lut (.A(n15008), .B(n14994), .C(\array[33] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2321[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_226_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_226_i5_3_lut_4_lut (.A(n15008), .B(n14994), .C(\array[33] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2321[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_226_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_226_i6_3_lut_4_lut (.A(n15008), .B(n14994), .C(\array[33] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2321[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_226_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_226_i7_3_lut_4_lut (.A(n15008), .B(n14994), .C(\array[33] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2321[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_226_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_226_i8_3_lut_4_lut (.A(n15008), .B(n14994), .C(\array[33] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2321[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_226_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_225_i1_3_lut_4_lut (.A(n15009), .B(n14994), .C(\array[34] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2329[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_225_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_225_i2_3_lut_4_lut (.A(n15009), .B(n14994), .C(\array[34] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2329[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_225_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_225_i3_3_lut_4_lut (.A(n15009), .B(n14994), .C(\array[34] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2329[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_225_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_225_i4_3_lut_4_lut (.A(n15009), .B(n14994), .C(\array[34] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2329[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_225_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_225_i5_3_lut_4_lut (.A(n15009), .B(n14994), .C(\array[34] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2329[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_225_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_225_i6_3_lut_4_lut (.A(n15009), .B(n14994), .C(\array[34] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2329[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_225_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_225_i7_3_lut_4_lut (.A(n15009), .B(n14994), .C(\array[34] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2329[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_225_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_225_i8_3_lut_4_lut (.A(n15009), .B(n14994), .C(\array[34] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2329[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_225_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_224_i1_3_lut_4_lut (.A(n15010), .B(n14994), .C(\array[35] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2337[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_224_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_224_i2_3_lut_4_lut (.A(n15010), .B(n14994), .C(\array[35] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2337[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_224_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_224_i3_3_lut_4_lut (.A(n15010), .B(n14994), .C(\array[35] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2337[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_224_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_224_i4_3_lut_4_lut (.A(n15010), .B(n14994), .C(\array[35] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2337[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_224_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_224_i5_3_lut_4_lut (.A(n15010), .B(n14994), .C(\array[35] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2337[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_224_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_224_i6_3_lut_4_lut (.A(n15010), .B(n14994), .C(\array[35] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2337[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_224_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_224_i7_3_lut_4_lut (.A(n15010), .B(n14994), .C(\array[35] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2337[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_224_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_224_i8_3_lut_4_lut (.A(n15010), .B(n14994), .C(\array[35] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2337[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_224_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_223_i1_3_lut_4_lut (.A(n15011), .B(n14994), .C(\array[36] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2345[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_223_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_223_i2_3_lut_4_lut (.A(n15011), .B(n14994), .C(\array[36] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2345[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_223_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_223_i3_3_lut_4_lut (.A(n15011), .B(n14994), .C(\array[36] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2345[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_223_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_223_i4_3_lut_4_lut (.A(n15011), .B(n14994), .C(\array[36] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2345[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_223_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_223_i5_3_lut_4_lut (.A(n15011), .B(n14994), .C(\array[36] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2345[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_223_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_223_i6_3_lut_4_lut (.A(n15011), .B(n14994), .C(\array[36] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2345[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_223_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_223_i7_3_lut_4_lut (.A(n15011), .B(n14994), .C(\array[36] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2345[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_223_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_223_i8_3_lut_4_lut (.A(n15011), .B(n14994), .C(\array[36] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2345[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_223_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_222_i1_3_lut_4_lut (.A(n15012), .B(n14994), .C(\array[37] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2353[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_222_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_222_i2_3_lut_4_lut (.A(n15012), .B(n14994), .C(\array[37] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2353[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_222_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_222_i3_3_lut_4_lut (.A(n15012), .B(n14994), .C(\array[37] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2353[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_222_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_222_i4_3_lut_4_lut (.A(n15012), .B(n14994), .C(\array[37] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2353[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_222_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_222_i5_3_lut_4_lut (.A(n15012), .B(n14994), .C(\array[37] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2353[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_222_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_222_i6_3_lut_4_lut (.A(n15012), .B(n14994), .C(\array[37] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2353[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_222_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_222_i7_3_lut_4_lut (.A(n15012), .B(n14994), .C(\array[37] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2353[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_222_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_222_i8_3_lut_4_lut (.A(n15012), .B(n14994), .C(\array[37] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2353[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_222_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_219_i1_3_lut_4_lut (.A(n15015), .B(n14994), .C(\array[40] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2377[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_219_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_219_i2_3_lut_4_lut (.A(n15015), .B(n14994), .C(\array[40] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2377[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_219_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_219_i3_3_lut_4_lut (.A(n15015), .B(n14994), .C(\array[40] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2377[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_219_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_219_i4_3_lut_4_lut (.A(n15015), .B(n14994), .C(\array[40] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2377[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_219_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_219_i5_3_lut_4_lut (.A(n15015), .B(n14994), .C(\array[40] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2377[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_219_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_219_i6_3_lut_4_lut (.A(n15015), .B(n14994), .C(\array[40] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2377[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_219_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_219_i7_3_lut_4_lut (.A(n15015), .B(n14994), .C(\array[40] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2377[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_219_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_219_i8_3_lut_4_lut (.A(n15015), .B(n14994), .C(\array[40] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2377[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_219_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_218_i1_3_lut_4_lut (.A(n15016), .B(n14994), .C(\array[41] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2385[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_218_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_218_i2_3_lut_4_lut (.A(n15016), .B(n14994), .C(\array[41] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2385[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_218_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_218_i3_3_lut_4_lut (.A(n15016), .B(n14994), .C(\array[41] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2385[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_218_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_218_i4_3_lut_4_lut (.A(n15016), .B(n14994), .C(\array[41] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2385[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_218_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_218_i5_3_lut_4_lut (.A(n15016), .B(n14994), .C(\array[41] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2385[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_218_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_218_i6_3_lut_4_lut (.A(n15016), .B(n14994), .C(\array[41] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2385[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_218_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_218_i7_3_lut_4_lut (.A(n15016), .B(n14994), .C(\array[41] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2385[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_218_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_218_i8_3_lut_4_lut (.A(n15016), .B(n14994), .C(\array[41] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2385[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_218_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_217_i1_3_lut_4_lut (.A(n15017), .B(n14994), .C(\array[42] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2393[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_217_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_217_i2_3_lut_4_lut (.A(n15017), .B(n14994), .C(\array[42] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2393[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_217_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_217_i3_3_lut_4_lut (.A(n15017), .B(n14994), .C(\array[42] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2393[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_217_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_217_i4_3_lut_4_lut (.A(n15017), .B(n14994), .C(\array[42] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2393[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_217_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_217_i5_3_lut_4_lut (.A(n15017), .B(n14994), .C(\array[42] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2393[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_217_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_217_i6_3_lut_4_lut (.A(n15017), .B(n14994), .C(\array[42] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2393[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_217_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_217_i7_3_lut_4_lut (.A(n15017), .B(n14994), .C(\array[42] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2393[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_217_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_217_i8_3_lut_4_lut (.A(n15017), .B(n14994), .C(\array[42] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2393[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_217_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_216_i1_3_lut_4_lut (.A(n15018), .B(n14994), .C(\array[43] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2401[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_216_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_216_i2_3_lut_4_lut (.A(n15018), .B(n14994), .C(\array[43] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2401[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_216_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_216_i3_3_lut_4_lut (.A(n15018), .B(n14994), .C(\array[43] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2401[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_216_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_216_i4_3_lut_4_lut (.A(n15018), .B(n14994), .C(\array[43] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2401[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_216_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_216_i5_3_lut_4_lut (.A(n15018), .B(n14994), .C(\array[43] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2401[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_216_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_216_i6_3_lut_4_lut (.A(n15018), .B(n14994), .C(\array[43] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2401[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_216_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_216_i7_3_lut_4_lut (.A(n15018), .B(n14994), .C(\array[43] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2401[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_216_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_216_i8_3_lut_4_lut (.A(n15018), .B(n14994), .C(\array[43] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2401[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_216_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_215_i1_3_lut_4_lut (.A(n15019), .B(n14994), .C(\array[44] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2409[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_215_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_215_i2_3_lut_4_lut (.A(n15019), .B(n14994), .C(\array[44] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2409[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_215_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_215_i3_3_lut_4_lut (.A(n15019), .B(n14994), .C(\array[44] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2409[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_215_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_215_i4_3_lut_4_lut (.A(n15019), .B(n14994), .C(\array[44] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2409[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_215_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_215_i5_3_lut_4_lut (.A(n15019), .B(n14994), .C(\array[44] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2409[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_215_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_215_i6_3_lut_4_lut (.A(n15019), .B(n14994), .C(\array[44] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2409[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_215_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_215_i7_3_lut_4_lut (.A(n15019), .B(n14994), .C(\array[44] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2409[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_215_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_215_i8_3_lut_4_lut (.A(n15019), .B(n14994), .C(\array[44] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2409[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_215_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_214_i1_3_lut_4_lut (.A(n15020), .B(n14994), .C(\array[45] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2417[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_214_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_214_i2_3_lut_4_lut (.A(n15020), .B(n14994), .C(\array[45] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2417[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_214_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_214_i3_3_lut_4_lut (.A(n15020), .B(n14994), .C(\array[45] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2417[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_214_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_214_i4_3_lut_4_lut (.A(n15020), .B(n14994), .C(\array[45] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2417[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_214_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_214_i5_3_lut_4_lut (.A(n15020), .B(n14994), .C(\array[45] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2417[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_214_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_214_i6_3_lut_4_lut (.A(n15020), .B(n14994), .C(\array[45] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2417[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_214_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_214_i7_3_lut_4_lut (.A(n15020), .B(n14994), .C(\array[45] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2417[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_214_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_214_i8_3_lut_4_lut (.A(n15020), .B(n14994), .C(\array[45] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2417[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_214_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_213_i1_3_lut_4_lut (.A(n15021), .B(n14994), .C(\array[46] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2425[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_213_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_213_i2_3_lut_4_lut (.A(n15021), .B(n14994), .C(\array[46] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2425[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_213_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_213_i3_3_lut_4_lut (.A(n15021), .B(n14994), .C(\array[46] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2425[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_213_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_213_i4_3_lut_4_lut (.A(n15021), .B(n14994), .C(\array[46] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2425[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_213_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_213_i5_3_lut_4_lut (.A(n15021), .B(n14994), .C(\array[46] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2425[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_213_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_213_i6_3_lut_4_lut (.A(n15021), .B(n14994), .C(\array[46] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2425[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_213_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_213_i7_3_lut_4_lut (.A(n15021), .B(n14994), .C(\array[46] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2425[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_213_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_213_i8_3_lut_4_lut (.A(n15021), .B(n14994), .C(\array[46] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2425[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_213_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_212_i1_3_lut_4_lut (.A(n15023), .B(n14994), .C(\array[47] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2433[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_212_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_212_i2_3_lut_4_lut (.A(n15023), .B(n14994), .C(\array[47] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2433[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_212_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_212_i3_3_lut_4_lut (.A(n15023), .B(n14994), .C(\array[47] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2433[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_212_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_212_i4_3_lut_4_lut (.A(n15023), .B(n14994), .C(\array[47] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2433[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_212_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_212_i5_3_lut_4_lut (.A(n15023), .B(n14994), .C(\array[47] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2433[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_212_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_212_i6_3_lut_4_lut (.A(n15023), .B(n14994), .C(\array[47] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2433[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_212_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_212_i7_3_lut_4_lut (.A(n15023), .B(n14994), .C(\array[47] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2433[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_212_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_212_i8_3_lut_4_lut (.A(n15023), .B(n14994), .C(\array[47] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2433[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_212_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_211_i1_3_lut_4_lut (.A(n15007), .B(n14995), .C(\array[48] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2441[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_211_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_211_i2_3_lut_4_lut (.A(n15007), .B(n14995), .C(\array[48] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2441[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_211_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_211_i3_3_lut_4_lut (.A(n15007), .B(n14995), .C(\array[48] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2441[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_211_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_211_i4_3_lut_4_lut (.A(n15007), .B(n14995), .C(\array[48] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2441[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_211_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_211_i5_3_lut_4_lut (.A(n15007), .B(n14995), .C(\array[48] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2441[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_211_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_211_i6_3_lut_4_lut (.A(n15007), .B(n14995), .C(\array[48] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2441[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_211_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_211_i7_3_lut_4_lut (.A(n15007), .B(n14995), .C(\array[48] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2441[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_211_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_211_i8_3_lut_4_lut (.A(n15007), .B(n14995), .C(\array[48] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2441[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_211_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_210_i1_3_lut_4_lut (.A(n15008), .B(n14995), .C(\array[49] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2449[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_210_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_210_i2_3_lut_4_lut (.A(n15008), .B(n14995), .C(\array[49] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2449[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_210_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_210_i3_3_lut_4_lut (.A(n15008), .B(n14995), .C(\array[49] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2449[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_210_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_210_i4_3_lut_4_lut (.A(n15008), .B(n14995), .C(\array[49] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2449[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_210_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_210_i5_3_lut_4_lut (.A(n15008), .B(n14995), .C(\array[49] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2449[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_210_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_210_i6_3_lut_4_lut (.A(n15008), .B(n14995), .C(\array[49] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2449[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_210_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_210_i7_3_lut_4_lut (.A(n15008), .B(n14995), .C(\array[49] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2449[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_210_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_210_i8_3_lut_4_lut (.A(n15008), .B(n14995), .C(\array[49] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2449[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_210_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_209_i1_3_lut_4_lut (.A(n15009), .B(n14995), .C(\array[50] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2457[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_209_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_209_i2_3_lut_4_lut (.A(n15009), .B(n14995), .C(\array[50] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2457[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_209_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_209_i3_3_lut_4_lut (.A(n15009), .B(n14995), .C(\array[50] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2457[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_209_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_209_i4_3_lut_4_lut (.A(n15009), .B(n14995), .C(\array[50] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2457[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_209_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_209_i5_3_lut_4_lut (.A(n15009), .B(n14995), .C(\array[50] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2457[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_209_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_209_i6_3_lut_4_lut (.A(n15009), .B(n14995), .C(\array[50] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2457[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_209_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_209_i7_3_lut_4_lut (.A(n15009), .B(n14995), .C(\array[50] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2457[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_209_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_209_i8_3_lut_4_lut (.A(n15009), .B(n14995), .C(\array[50] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2457[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_209_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_208_i1_3_lut_4_lut (.A(n15010), .B(n14995), .C(\array[51] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2465[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_208_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_208_i2_3_lut_4_lut (.A(n15010), .B(n14995), .C(\array[51] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2465[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_208_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_208_i3_3_lut_4_lut (.A(n15010), .B(n14995), .C(\array[51] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2465[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_208_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_208_i4_3_lut_4_lut (.A(n15010), .B(n14995), .C(\array[51] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2465[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_208_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_208_i5_3_lut_4_lut (.A(n15010), .B(n14995), .C(\array[51] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2465[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_208_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_208_i6_3_lut_4_lut (.A(n15010), .B(n14995), .C(\array[51] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2465[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_208_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_208_i7_3_lut_4_lut (.A(n15010), .B(n14995), .C(\array[51] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2465[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_208_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_208_i8_3_lut_4_lut (.A(n15010), .B(n14995), .C(\array[51] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2465[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_208_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_207_i1_3_lut_4_lut (.A(n15011), .B(n14995), .C(\array[52] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2473[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_207_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_207_i2_3_lut_4_lut (.A(n15011), .B(n14995), .C(\array[52] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2473[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_207_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_207_i3_3_lut_4_lut (.A(n15011), .B(n14995), .C(\array[52] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2473[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_207_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_207_i4_3_lut_4_lut (.A(n15011), .B(n14995), .C(\array[52] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2473[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_207_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_207_i5_3_lut_4_lut (.A(n15011), .B(n14995), .C(\array[52] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2473[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_207_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_207_i6_3_lut_4_lut (.A(n15011), .B(n14995), .C(\array[52] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2473[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_207_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_207_i7_3_lut_4_lut (.A(n15011), .B(n14995), .C(\array[52] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2473[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_207_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_207_i8_3_lut_4_lut (.A(n15011), .B(n14995), .C(\array[52] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2473[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_207_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_206_i1_3_lut_4_lut (.A(n15012), .B(n14995), .C(\array[53] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2481[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_206_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_206_i2_3_lut_4_lut (.A(n15012), .B(n14995), .C(\array[53] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2481[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_206_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_206_i3_3_lut_4_lut (.A(n15012), .B(n14995), .C(\array[53] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2481[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_206_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_206_i4_3_lut_4_lut (.A(n15012), .B(n14995), .C(\array[53] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2481[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_206_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_206_i5_3_lut_4_lut (.A(n15012), .B(n14995), .C(\array[53] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2481[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_206_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_206_i6_3_lut_4_lut (.A(n15012), .B(n14995), .C(\array[53] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2481[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_206_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_206_i7_3_lut_4_lut (.A(n15012), .B(n14995), .C(\array[53] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2481[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_206_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_206_i8_3_lut_4_lut (.A(n15012), .B(n14995), .C(\array[53] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2481[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_206_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_205_i1_3_lut_4_lut (.A(n15013), .B(n14995), .C(\array[54] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2489[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_205_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_205_i2_3_lut_4_lut (.A(n15013), .B(n14995), .C(\array[54] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2489[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_205_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_205_i3_3_lut_4_lut (.A(n15013), .B(n14995), .C(\array[54] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2489[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_205_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_205_i4_3_lut_4_lut (.A(n15013), .B(n14995), .C(\array[54] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2489[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_205_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_205_i5_3_lut_4_lut (.A(n15013), .B(n14995), .C(\array[54] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2489[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_205_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_205_i6_3_lut_4_lut (.A(n15013), .B(n14995), .C(\array[54] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2489[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_205_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_205_i7_3_lut_4_lut (.A(n15013), .B(n14995), .C(\array[54] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2489[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_205_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_205_i8_3_lut_4_lut (.A(n15013), .B(n14995), .C(\array[54] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2489[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_205_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_204_i1_3_lut_4_lut (.A(n15014), .B(n14995), .C(\array[55] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2497[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_204_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_204_i2_3_lut_4_lut (.A(n15014), .B(n14995), .C(\array[55] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2497[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_204_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_204_i3_3_lut_4_lut (.A(n15014), .B(n14995), .C(\array[55] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2497[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_204_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_204_i4_3_lut_4_lut (.A(n15014), .B(n14995), .C(\array[55] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2497[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_204_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_204_i5_3_lut_4_lut (.A(n15014), .B(n14995), .C(\array[55] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2497[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_204_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_204_i6_3_lut_4_lut (.A(n15014), .B(n14995), .C(\array[55] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2497[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_204_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_204_i7_3_lut_4_lut (.A(n15014), .B(n14995), .C(\array[55] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2497[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_204_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_204_i8_3_lut_4_lut (.A(n15014), .B(n14995), .C(\array[55] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2497[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_204_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_203_i1_3_lut_4_lut (.A(n15015), .B(n14995), .C(\array[56] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2505[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_203_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_203_i2_3_lut_4_lut (.A(n15015), .B(n14995), .C(\array[56] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2505[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_203_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_203_i3_3_lut_4_lut (.A(n15015), .B(n14995), .C(\array[56] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2505[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_203_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_203_i4_3_lut_4_lut (.A(n15015), .B(n14995), .C(\array[56] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2505[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_203_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_203_i5_3_lut_4_lut (.A(n15015), .B(n14995), .C(\array[56] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2505[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_203_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_203_i6_3_lut_4_lut (.A(n15015), .B(n14995), .C(\array[56] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2505[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_203_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_203_i7_3_lut_4_lut (.A(n15015), .B(n14995), .C(\array[56] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2505[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_203_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_203_i8_3_lut_4_lut (.A(n15015), .B(n14995), .C(\array[56] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2505[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_203_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_202_i1_3_lut_4_lut (.A(n15016), .B(n14995), .C(\array[57] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2513[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_202_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_202_i2_3_lut_4_lut (.A(n15016), .B(n14995), .C(\array[57] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2513[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_202_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_202_i3_3_lut_4_lut (.A(n15016), .B(n14995), .C(\array[57] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2513[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_202_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_202_i4_3_lut_4_lut (.A(n15016), .B(n14995), .C(\array[57] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2513[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_202_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_202_i5_3_lut_4_lut (.A(n15016), .B(n14995), .C(\array[57] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2513[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_202_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_202_i6_3_lut_4_lut (.A(n15016), .B(n14995), .C(\array[57] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2513[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_202_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_202_i7_3_lut_4_lut (.A(n15016), .B(n14995), .C(\array[57] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2513[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_202_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_202_i8_3_lut_4_lut (.A(n15016), .B(n14995), .C(\array[57] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2513[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_202_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_201_i1_3_lut_4_lut (.A(n15017), .B(n14995), .C(\array[58] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2521[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_201_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_201_i2_3_lut_4_lut (.A(n15017), .B(n14995), .C(\array[58] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2521[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_201_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_201_i3_3_lut_4_lut (.A(n15017), .B(n14995), .C(\array[58] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2521[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_201_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_201_i4_3_lut_4_lut (.A(n15017), .B(n14995), .C(\array[58] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2521[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_201_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_201_i5_3_lut_4_lut (.A(n15017), .B(n14995), .C(\array[58] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2521[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_201_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_201_i6_3_lut_4_lut (.A(n15017), .B(n14995), .C(\array[58] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2521[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_201_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_201_i7_3_lut_4_lut (.A(n15017), .B(n14995), .C(\array[58] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2521[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_201_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_201_i8_3_lut_4_lut (.A(n15017), .B(n14995), .C(\array[58] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2521[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_201_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_200_i1_3_lut_4_lut (.A(n15018), .B(n14995), .C(\array[59] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2529[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_200_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_200_i2_3_lut_4_lut (.A(n15018), .B(n14995), .C(\array[59] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2529[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_200_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_200_i3_3_lut_4_lut (.A(n15018), .B(n14995), .C(\array[59] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2529[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_200_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_200_i4_3_lut_4_lut (.A(n15018), .B(n14995), .C(\array[59] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2529[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_200_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_200_i5_3_lut_4_lut (.A(n15018), .B(n14995), .C(\array[59] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2529[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_200_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_200_i6_3_lut_4_lut (.A(n15018), .B(n14995), .C(\array[59] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2529[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_200_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_200_i7_3_lut_4_lut (.A(n15018), .B(n14995), .C(\array[59] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2529[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_200_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_200_i8_3_lut_4_lut (.A(n15018), .B(n14995), .C(\array[59] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2529[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_200_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_199_i1_3_lut_4_lut (.A(n15019), .B(n14995), .C(\array[60] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2537[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_199_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_199_i2_3_lut_4_lut (.A(n15019), .B(n14995), .C(\array[60] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2537[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_199_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_199_i3_3_lut_4_lut (.A(n15019), .B(n14995), .C(\array[60] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2537[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_199_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_199_i4_3_lut_4_lut (.A(n15019), .B(n14995), .C(\array[60] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2537[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_199_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_199_i5_3_lut_4_lut (.A(n15019), .B(n14995), .C(\array[60] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2537[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_199_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_199_i6_3_lut_4_lut (.A(n15019), .B(n14995), .C(\array[60] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2537[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_199_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_199_i7_3_lut_4_lut (.A(n15019), .B(n14995), .C(\array[60] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2537[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_199_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_199_i8_3_lut_4_lut (.A(n15019), .B(n14995), .C(\array[60] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2537[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_199_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_198_i1_3_lut_4_lut (.A(n15020), .B(n14995), .C(\array[61] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2545[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_198_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_198_i2_3_lut_4_lut (.A(n15020), .B(n14995), .C(\array[61] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2545[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_198_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_198_i3_3_lut_4_lut (.A(n15020), .B(n14995), .C(\array[61] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2545[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_198_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_198_i4_3_lut_4_lut (.A(n15020), .B(n14995), .C(\array[61] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2545[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_198_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_198_i5_3_lut_4_lut (.A(n15020), .B(n14995), .C(\array[61] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2545[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_198_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_198_i6_3_lut_4_lut (.A(n15020), .B(n14995), .C(\array[61] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2545[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_198_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_198_i7_3_lut_4_lut (.A(n15020), .B(n14995), .C(\array[61] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2545[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_198_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_198_i8_3_lut_4_lut (.A(n15020), .B(n14995), .C(\array[61] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2545[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_198_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_197_i1_3_lut_4_lut (.A(n15021), .B(n14995), .C(\array[62] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2553[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_197_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_197_i2_3_lut_4_lut (.A(n15021), .B(n14995), .C(\array[62] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2553[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_197_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_197_i3_3_lut_4_lut (.A(n15021), .B(n14995), .C(\array[62] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2553[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_197_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_197_i4_3_lut_4_lut (.A(n15021), .B(n14995), .C(\array[62] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2553[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_197_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_197_i5_3_lut_4_lut (.A(n15021), .B(n14995), .C(\array[62] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2553[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_197_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_197_i6_3_lut_4_lut (.A(n15021), .B(n14995), .C(\array[62] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2553[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_197_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_197_i7_3_lut_4_lut (.A(n15021), .B(n14995), .C(\array[62] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2553[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_197_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_197_i8_3_lut_4_lut (.A(n15021), .B(n14995), .C(\array[62] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2553[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_197_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_196_i1_3_lut_4_lut (.A(n15023), .B(n14995), .C(\array[63] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2561[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_196_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_196_i2_3_lut_4_lut (.A(n15023), .B(n14995), .C(\array[63] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2561[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_196_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_196_i3_3_lut_4_lut (.A(n15023), .B(n14995), .C(\array[63] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2561[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_196_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_196_i4_3_lut_4_lut (.A(n15023), .B(n14995), .C(\array[63] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2561[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_196_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_196_i5_3_lut_4_lut (.A(n15023), .B(n14995), .C(\array[63] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2561[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_196_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_196_i6_3_lut_4_lut (.A(n15023), .B(n14995), .C(\array[63] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2561[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_196_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_196_i7_3_lut_4_lut (.A(n15023), .B(n14995), .C(\array[63] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2561[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_196_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_196_i8_3_lut_4_lut (.A(n15023), .B(n14995), .C(\array[63] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2561[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_196_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_195_i1_3_lut_4_lut (.A(n15007), .B(n14996), .C(\array[64] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2569[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_195_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_195_i2_3_lut_4_lut (.A(n15007), .B(n14996), .C(\array[64] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2569[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_195_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_195_i3_3_lut_4_lut (.A(n15007), .B(n14996), .C(\array[64] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2569[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_195_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_195_i4_3_lut_4_lut (.A(n15007), .B(n14996), .C(\array[64] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2569[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_195_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_195_i5_3_lut_4_lut (.A(n15007), .B(n14996), .C(\array[64] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2569[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_195_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_195_i6_3_lut_4_lut (.A(n15007), .B(n14996), .C(\array[64] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2569[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_195_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_195_i7_3_lut_4_lut (.A(n15007), .B(n14996), .C(\array[64] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2569[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_195_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_195_i8_3_lut_4_lut (.A(n15007), .B(n14996), .C(\array[64] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2569[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_195_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_194_i1_3_lut_4_lut (.A(n15008), .B(n14996), .C(\array[65] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2577[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_194_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_194_i2_3_lut_4_lut (.A(n15008), .B(n14996), .C(\array[65] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2577[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_194_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_194_i3_3_lut_4_lut (.A(n15008), .B(n14996), .C(\array[65] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2577[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_194_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_194_i4_3_lut_4_lut (.A(n15008), .B(n14996), .C(\array[65] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2577[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_194_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_194_i5_3_lut_4_lut (.A(n15008), .B(n14996), .C(\array[65] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2577[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_194_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_194_i6_3_lut_4_lut (.A(n15008), .B(n14996), .C(\array[65] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2577[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_194_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_194_i7_3_lut_4_lut (.A(n15008), .B(n14996), .C(\array[65] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2577[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_194_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_194_i8_3_lut_4_lut (.A(n15008), .B(n14996), .C(\array[65] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2577[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_194_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_193_i1_3_lut_4_lut (.A(n15009), .B(n14996), .C(\array[66] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2585[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_193_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_193_i2_3_lut_4_lut (.A(n15009), .B(n14996), .C(\array[66] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2585[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_193_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_193_i3_3_lut_4_lut (.A(n15009), .B(n14996), .C(\array[66] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2585[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_193_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_193_i4_3_lut_4_lut (.A(n15009), .B(n14996), .C(\array[66] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2585[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_193_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_193_i5_3_lut_4_lut (.A(n15009), .B(n14996), .C(\array[66] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2585[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_193_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_193_i6_3_lut_4_lut (.A(n15009), .B(n14996), .C(\array[66] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2585[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_193_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_193_i7_3_lut_4_lut (.A(n15009), .B(n14996), .C(\array[66] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2585[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_193_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_193_i8_3_lut_4_lut (.A(n15009), .B(n14996), .C(\array[66] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2585[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_193_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_192_i1_3_lut_4_lut (.A(n15010), .B(n14996), .C(\array[67] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2593[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_192_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_192_i2_3_lut_4_lut (.A(n15010), .B(n14996), .C(\array[67] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2593[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_192_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_192_i3_3_lut_4_lut (.A(n15010), .B(n14996), .C(\array[67] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2593[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_192_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_192_i4_3_lut_4_lut (.A(n15010), .B(n14996), .C(\array[67] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2593[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_192_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_192_i5_3_lut_4_lut (.A(n15010), .B(n14996), .C(\array[67] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2593[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_192_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_192_i6_3_lut_4_lut (.A(n15010), .B(n14996), .C(\array[67] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2593[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_192_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_192_i7_3_lut_4_lut (.A(n15010), .B(n14996), .C(\array[67] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2593[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_192_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_192_i8_3_lut_4_lut (.A(n15010), .B(n14996), .C(\array[67] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2593[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_192_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_191_i1_3_lut_4_lut (.A(n15011), .B(n14996), .C(\array[68] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2601[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_191_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_191_i2_3_lut_4_lut (.A(n15011), .B(n14996), .C(\array[68] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2601[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_191_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_191_i3_3_lut_4_lut (.A(n15011), .B(n14996), .C(\array[68] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2601[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_191_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_191_i4_3_lut_4_lut (.A(n15011), .B(n14996), .C(\array[68] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2601[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_191_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_191_i5_3_lut_4_lut (.A(n15011), .B(n14996), .C(\array[68] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2601[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_191_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_191_i6_3_lut_4_lut (.A(n15011), .B(n14996), .C(\array[68] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2601[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_191_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_191_i7_3_lut_4_lut (.A(n15011), .B(n14996), .C(\array[68] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2601[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_191_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_191_i8_3_lut_4_lut (.A(n15011), .B(n14996), .C(\array[68] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2601[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_191_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_190_i1_3_lut_4_lut (.A(n15012), .B(n14996), .C(\array[69] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2609[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_190_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_190_i2_3_lut_4_lut (.A(n15012), .B(n14996), .C(\array[69] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2609[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_190_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_190_i3_3_lut_4_lut (.A(n15012), .B(n14996), .C(\array[69] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2609[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_190_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_190_i4_3_lut_4_lut (.A(n15012), .B(n14996), .C(\array[69] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2609[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_190_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_190_i5_3_lut_4_lut (.A(n15012), .B(n14996), .C(\array[69] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2609[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_190_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_190_i6_3_lut_4_lut (.A(n15012), .B(n14996), .C(\array[69] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2609[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_190_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_190_i7_3_lut_4_lut (.A(n15012), .B(n14996), .C(\array[69] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2609[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_190_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_190_i8_3_lut_4_lut (.A(n15012), .B(n14996), .C(\array[69] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2609[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_190_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_189_i1_3_lut_4_lut (.A(n15013), .B(n14996), .C(\array[70] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2617[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_189_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_189_i2_3_lut_4_lut (.A(n15013), .B(n14996), .C(\array[70] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2617[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_189_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_189_i3_3_lut_4_lut (.A(n15013), .B(n14996), .C(\array[70] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2617[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_189_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_189_i4_3_lut_4_lut (.A(n15013), .B(n14996), .C(\array[70] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2617[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_189_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_189_i5_3_lut_4_lut (.A(n15013), .B(n14996), .C(\array[70] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2617[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_189_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_189_i6_3_lut_4_lut (.A(n15013), .B(n14996), .C(\array[70] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2617[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_189_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_189_i7_3_lut_4_lut (.A(n15013), .B(n14996), .C(\array[70] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2617[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_189_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_189_i8_3_lut_4_lut (.A(n15013), .B(n14996), .C(\array[70] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2617[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_189_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_188_i1_3_lut_4_lut (.A(n15014), .B(n14996), .C(\array[71] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2625[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_188_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_188_i2_3_lut_4_lut (.A(n15014), .B(n14996), .C(\array[71] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2625[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_188_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_188_i3_3_lut_4_lut (.A(n15014), .B(n14996), .C(\array[71] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2625[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_188_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_188_i4_3_lut_4_lut (.A(n15014), .B(n14996), .C(\array[71] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2625[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_188_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_188_i5_3_lut_4_lut (.A(n15014), .B(n14996), .C(\array[71] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2625[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_188_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_188_i6_3_lut_4_lut (.A(n15014), .B(n14996), .C(\array[71] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2625[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_188_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_188_i7_3_lut_4_lut (.A(n15014), .B(n14996), .C(\array[71] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2625[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_188_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_188_i8_3_lut_4_lut (.A(n15014), .B(n14996), .C(\array[71] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2625[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_188_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_187_i1_3_lut_4_lut (.A(n15015), .B(n14996), .C(\array[72] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2633[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_187_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_187_i2_3_lut_4_lut (.A(n15015), .B(n14996), .C(\array[72] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2633[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_187_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_187_i3_3_lut_4_lut (.A(n15015), .B(n14996), .C(\array[72] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2633[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_187_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_187_i4_3_lut_4_lut (.A(n15015), .B(n14996), .C(\array[72] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2633[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_187_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_187_i5_3_lut_4_lut (.A(n15015), .B(n14996), .C(\array[72] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2633[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_187_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_187_i6_3_lut_4_lut (.A(n15015), .B(n14996), .C(\array[72] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2633[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_187_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_187_i7_3_lut_4_lut (.A(n15015), .B(n14996), .C(\array[72] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2633[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_187_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_187_i8_3_lut_4_lut (.A(n15015), .B(n14996), .C(\array[72] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2633[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_187_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_186_i1_3_lut_4_lut (.A(n15016), .B(n14996), .C(\array[73] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2641[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_186_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_186_i2_3_lut_4_lut (.A(n15016), .B(n14996), .C(\array[73] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2641[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_186_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 wr_en_pad_lut_buf_2 (.A(wr_en_c), .Z(clk_c_enable_2007)) /* synthesis lut_function=(A) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(17[16:21])
    defparam wr_en_pad_lut_buf_2.init = 16'haaaa;
    LUT4 mux_186_i3_3_lut_4_lut (.A(n15016), .B(n14996), .C(\array[73] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2641[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_186_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_186_i4_3_lut_4_lut (.A(n15016), .B(n14996), .C(\array[73] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2641[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_186_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_186_i5_3_lut_4_lut (.A(n15016), .B(n14996), .C(\array[73] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2641[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_186_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_186_i6_3_lut_4_lut (.A(n15016), .B(n14996), .C(\array[73] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2641[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_186_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 wr_en_pad_lut_buf_1 (.A(wr_en_c), .Z(clk_c_enable_1007)) /* synthesis lut_function=(A) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(17[16:21])
    defparam wr_en_pad_lut_buf_1.init = 16'haaaa;
    LUT4 mux_186_i7_3_lut_4_lut (.A(n15016), .B(n14996), .C(\array[73] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2641[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_186_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_186_i8_3_lut_4_lut (.A(n15016), .B(n14996), .C(\array[73] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2641[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_186_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_185_i1_3_lut_4_lut (.A(n15017), .B(n14996), .C(\array[74] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2649[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_185_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_185_i2_3_lut_4_lut (.A(n15017), .B(n14996), .C(\array[74] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2649[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_185_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_185_i3_3_lut_4_lut (.A(n15017), .B(n14996), .C(\array[74] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2649[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_185_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_185_i4_3_lut_4_lut (.A(n15017), .B(n14996), .C(\array[74] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2649[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_185_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_185_i5_3_lut_4_lut (.A(n15017), .B(n14996), .C(\array[74] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2649[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_185_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 wr_en_pad_lut_buf_3 (.A(wr_en_c), .Z(clk_c_enable_2056)) /* synthesis lut_function=(A) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(17[16:21])
    defparam wr_en_pad_lut_buf_3.init = 16'haaaa;
    LUT4 mux_185_i6_3_lut_4_lut (.A(n15017), .B(n14996), .C(\array[74] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2649[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_185_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_185_i7_3_lut_4_lut (.A(n15017), .B(n14996), .C(\array[74] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2649[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_185_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_185_i8_3_lut_4_lut (.A(n15017), .B(n14996), .C(\array[74] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2649[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_185_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_184_i1_3_lut_4_lut (.A(n15018), .B(n14996), .C(\array[75] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2657[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_184_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_184_i2_3_lut_4_lut (.A(n15018), .B(n14996), .C(\array[75] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2657[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_184_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_184_i3_3_lut_4_lut (.A(n15018), .B(n14996), .C(\array[75] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2657[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_184_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_184_i4_3_lut_4_lut (.A(n15018), .B(n14996), .C(\array[75] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2657[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_184_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_184_i5_3_lut_4_lut (.A(n15018), .B(n14996), .C(\array[75] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2657[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_184_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_184_i6_3_lut_4_lut (.A(n15018), .B(n14996), .C(\array[75] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2657[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_184_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_184_i7_3_lut_4_lut (.A(n15018), .B(n14996), .C(\array[75] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2657[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_184_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_184_i8_3_lut_4_lut (.A(n15018), .B(n14996), .C(\array[75] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2657[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_184_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_183_i1_3_lut_4_lut (.A(n15019), .B(n14996), .C(\array[76] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2665[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_183_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_183_i2_3_lut_4_lut (.A(n15019), .B(n14996), .C(\array[76] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2665[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_183_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_183_i3_3_lut_4_lut (.A(n15019), .B(n14996), .C(\array[76] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2665[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_183_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_183_i4_3_lut_4_lut (.A(n15019), .B(n14996), .C(\array[76] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2665[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_183_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_183_i5_3_lut_4_lut (.A(n15019), .B(n14996), .C(\array[76] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2665[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_183_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_511_i14_2_lut_rep_44_3_lut_4_lut (.A(addr_c_4), .B(addr_c_5), 
         .C(addr_c_7), .D(addr_c_6), .Z(n14992)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_511_i14_2_lut_rep_44_3_lut_4_lut.init = 16'hfffe;
    LUT4 equal_447_i14_2_lut_rep_48_3_lut_4_lut (.A(addr_c_4), .B(addr_c_5), 
         .C(addr_c_7), .D(addr_c_6), .Z(n14996)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_447_i14_2_lut_rep_48_3_lut_4_lut.init = 16'hfeff;
    LUT4 equal_383_i14_2_lut_rep_52_3_lut_4_lut (.A(addr_c_4), .B(addr_c_5), 
         .C(addr_c_7), .D(addr_c_6), .Z(n15000)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_383_i14_2_lut_rep_52_3_lut_4_lut.init = 16'hffef;
    LUT4 mux_183_i6_3_lut_4_lut (.A(n15019), .B(n14996), .C(\array[76] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2665[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_183_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_183_i7_3_lut_4_lut (.A(n15019), .B(n14996), .C(\array[76] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2665[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_183_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_183_i8_3_lut_4_lut (.A(n15019), .B(n14996), .C(\array[76] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2665[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_183_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_182_i1_3_lut_4_lut (.A(n15020), .B(n14996), .C(\array[77] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2673[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_182_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_182_i2_3_lut_4_lut (.A(n15020), .B(n14996), .C(\array[77] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2673[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_182_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_182_i3_3_lut_4_lut (.A(n15020), .B(n14996), .C(\array[77] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2673[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_182_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_182_i4_3_lut_4_lut (.A(n15020), .B(n14996), .C(\array[77] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2673[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_182_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_495_i14_2_lut_rep_45_3_lut_4_lut (.A(addr_c_4), .B(addr_c_5), 
         .C(addr_c_7), .D(addr_c_6), .Z(n14993)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_495_i14_2_lut_rep_45_3_lut_4_lut.init = 16'hfffd;
    LUT4 equal_367_i14_2_lut_rep_53_3_lut_4_lut (.A(addr_c_4), .B(addr_c_5), 
         .C(addr_c_7), .D(addr_c_6), .Z(n15001)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_367_i14_2_lut_rep_53_3_lut_4_lut.init = 16'hffdf;
    LUT4 mux_182_i5_3_lut_4_lut (.A(n15020), .B(n14996), .C(\array[77] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2673[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_182_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_431_i14_2_lut_rep_49_3_lut_4_lut (.A(addr_c_4), .B(addr_c_5), 
         .C(addr_c_7), .D(addr_c_6), .Z(n14997)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_431_i14_2_lut_rep_49_3_lut_4_lut.init = 16'hfdff;
    LUT4 mux_182_i6_3_lut_4_lut (.A(n15020), .B(n14996), .C(\array[77] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2673[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_182_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_182_i7_3_lut_4_lut (.A(n15020), .B(n14996), .C(\array[77] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2673[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_182_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_182_i8_3_lut_4_lut (.A(n15020), .B(n14996), .C(\array[77] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2673[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_182_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_181_i1_3_lut_4_lut (.A(n15021), .B(n14996), .C(\array[78] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2681[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_181_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_181_i2_3_lut_4_lut (.A(n15021), .B(n14996), .C(\array[78] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2681[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_181_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_479_i14_2_lut_rep_46_3_lut_4_lut (.A(addr_c_4), .B(addr_c_5), 
         .C(addr_c_7), .D(addr_c_6), .Z(n14994)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_479_i14_2_lut_rep_46_3_lut_4_lut.init = 16'hfffb;
    LUT4 equal_415_i14_2_lut_rep_50_3_lut_4_lut (.A(addr_c_4), .B(addr_c_5), 
         .C(addr_c_7), .D(addr_c_6), .Z(n14998)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_415_i14_2_lut_rep_50_3_lut_4_lut.init = 16'hfbff;
    LUT4 mux_181_i3_3_lut_4_lut (.A(n15021), .B(n14996), .C(\array[78] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2681[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_181_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_181_i4_3_lut_4_lut (.A(n15021), .B(n14996), .C(\array[78] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2681[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_181_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_181_i5_3_lut_4_lut (.A(n15021), .B(n14996), .C(\array[78] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2681[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_181_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_181_i6_3_lut_4_lut (.A(n15021), .B(n14996), .C(\array[78] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2681[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_181_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_181_i7_3_lut_4_lut (.A(n15021), .B(n14996), .C(\array[78] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2681[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_181_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_351_i14_2_lut_rep_54_3_lut_4_lut (.A(addr_c_4), .B(addr_c_5), 
         .C(addr_c_7), .D(addr_c_6), .Z(n15002)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_351_i14_2_lut_rep_54_3_lut_4_lut.init = 16'hffbf;
    LUT4 mux_181_i8_3_lut_4_lut (.A(n15021), .B(n14996), .C(\array[78] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2681[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_181_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_180_i1_3_lut_4_lut (.A(n15023), .B(n14996), .C(\array[79] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2689[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_180_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_180_i2_3_lut_4_lut (.A(n15023), .B(n14996), .C(\array[79] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2689[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_180_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_180_i3_3_lut_4_lut (.A(n15023), .B(n14996), .C(\array[79] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2689[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_180_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_180_i4_3_lut_4_lut (.A(n15023), .B(n14996), .C(\array[79] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2689[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_180_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_180_i5_3_lut_4_lut (.A(n15023), .B(n14996), .C(\array[79] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2689[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_180_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_180_i6_3_lut_4_lut (.A(n15023), .B(n14996), .C(\array[79] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2689[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_180_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_180_i7_3_lut_4_lut (.A(n15023), .B(n14996), .C(\array[79] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2689[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_180_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_180_i8_3_lut_4_lut (.A(n15023), .B(n14996), .C(\array[79] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2689[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_180_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_179_i1_3_lut_4_lut (.A(n15007), .B(n14997), .C(\array[80] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2697[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_179_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_179_i2_3_lut_4_lut (.A(n15007), .B(n14997), .C(\array[80] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2697[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_179_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_179_i3_3_lut_4_lut (.A(n15007), .B(n14997), .C(\array[80] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2697[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_179_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_179_i4_3_lut_4_lut (.A(n15007), .B(n14997), .C(\array[80] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2697[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_179_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_179_i5_3_lut_4_lut (.A(n15007), .B(n14997), .C(\array[80] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2697[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_179_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_179_i6_3_lut_4_lut (.A(n15007), .B(n14997), .C(\array[80] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2697[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_179_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_179_i7_3_lut_4_lut (.A(n15007), .B(n14997), .C(\array[80] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2697[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_179_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_179_i8_3_lut_4_lut (.A(n15007), .B(n14997), .C(\array[80] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2697[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_179_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_178_i1_3_lut_4_lut (.A(n15008), .B(n14997), .C(\array[81] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2705[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_178_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_178_i2_3_lut_4_lut (.A(n15008), .B(n14997), .C(\array[81] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2705[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_178_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_178_i3_3_lut_4_lut (.A(n15008), .B(n14997), .C(\array[81] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2705[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_178_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_178_i4_3_lut_4_lut (.A(n15008), .B(n14997), .C(\array[81] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2705[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_178_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_178_i5_3_lut_4_lut (.A(n15008), .B(n14997), .C(\array[81] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2705[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_178_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_178_i6_3_lut_4_lut (.A(n15008), .B(n14997), .C(\array[81] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2705[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_178_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_278_i11_2_lut_rep_67_3_lut_4_lut (.A(addr_c_0), .B(addr_c_1), 
         .C(addr_c_3), .D(addr_c_2), .Z(n15015)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_278_i11_2_lut_rep_67_3_lut_4_lut.init = 16'hffef;
    LUT4 mux_178_i7_3_lut_4_lut (.A(n15008), .B(n14997), .C(\array[81] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2705[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_178_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_178_i8_3_lut_4_lut (.A(n15008), .B(n14997), .C(\array[81] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2705[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_178_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_286_i11_2_lut_rep_59_3_lut_4_lut (.A(addr_c_0), .B(addr_c_1), 
         .C(addr_c_3), .D(addr_c_2), .Z(n15007)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_286_i11_2_lut_rep_59_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_177_i1_3_lut_4_lut (.A(n15009), .B(n14997), .C(\array[82] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2713[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_177_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_177_i2_3_lut_4_lut (.A(n15009), .B(n14997), .C(\array[82] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2713[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_177_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_177_i3_3_lut_4_lut (.A(n15009), .B(n14997), .C(\array[82] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2713[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_177_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_282_i11_2_lut_rep_63_3_lut_4_lut (.A(addr_c_0), .B(addr_c_1), 
         .C(addr_c_3), .D(addr_c_2), .Z(n15011)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_282_i11_2_lut_rep_63_3_lut_4_lut.init = 16'hfeff;
    LUT4 mux_177_i4_3_lut_4_lut (.A(n15009), .B(n14997), .C(\array[82] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2713[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_177_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_177_i5_3_lut_4_lut (.A(n15009), .B(n14997), .C(\array[82] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2713[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_177_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_177_i6_3_lut_4_lut (.A(n15009), .B(n14997), .C(\array[82] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2713[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_177_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_177_i7_3_lut_4_lut (.A(n15009), .B(n14997), .C(\array[82] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2713[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_177_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_277_i11_2_lut_rep_68_3_lut_4_lut (.A(addr_c_0), .B(addr_c_1), 
         .C(addr_c_3), .D(addr_c_2), .Z(n15016)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_277_i11_2_lut_rep_68_3_lut_4_lut.init = 16'hffdf;
    LUT4 mux_177_i8_3_lut_4_lut (.A(n15009), .B(n14997), .C(\array[82] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2713[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_177_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_176_i1_3_lut_4_lut (.A(n15010), .B(n14997), .C(\array[83] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2721[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_176_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_176_i2_3_lut_4_lut (.A(n15010), .B(n14997), .C(\array[83] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2721[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_176_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_285_i11_2_lut_rep_60_3_lut_4_lut (.A(addr_c_0), .B(addr_c_1), 
         .C(addr_c_3), .D(addr_c_2), .Z(n15008)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_285_i11_2_lut_rep_60_3_lut_4_lut.init = 16'hfffd;
    LUT4 equal_281_i11_2_lut_rep_64_3_lut_4_lut (.A(addr_c_0), .B(addr_c_1), 
         .C(addr_c_3), .D(addr_c_2), .Z(n15012)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_281_i11_2_lut_rep_64_3_lut_4_lut.init = 16'hfdff;
    LUT4 equal_284_i11_2_lut_rep_61_3_lut_4_lut (.A(addr_c_0), .B(addr_c_1), 
         .C(addr_c_3), .D(addr_c_2), .Z(n15009)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_284_i11_2_lut_rep_61_3_lut_4_lut.init = 16'hfffb;
    LUT4 equal_276_i11_2_lut_rep_69_3_lut_4_lut (.A(addr_c_0), .B(addr_c_1), 
         .C(addr_c_3), .D(addr_c_2), .Z(n15017)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_276_i11_2_lut_rep_69_3_lut_4_lut.init = 16'hffbf;
    LUT4 mux_176_i3_3_lut_4_lut (.A(n15010), .B(n14997), .C(\array[83] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2721[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_176_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_176_i4_3_lut_4_lut (.A(n15010), .B(n14997), .C(\array[83] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2721[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_176_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_176_i5_3_lut_4_lut (.A(n15010), .B(n14997), .C(\array[83] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2721[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_176_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_176_i6_3_lut_4_lut (.A(n15010), .B(n14997), .C(\array[83] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2721[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_176_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_176_i7_3_lut_4_lut (.A(n15010), .B(n14997), .C(\array[83] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2721[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_176_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_176_i8_3_lut_4_lut (.A(n15010), .B(n14997), .C(\array[83] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2721[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_176_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_280_i11_2_lut_rep_65_3_lut_4_lut (.A(addr_c_0), .B(addr_c_1), 
         .C(addr_c_3), .D(addr_c_2), .Z(n15013)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam equal_280_i11_2_lut_rep_65_3_lut_4_lut.init = 16'hfbff;
    LUT4 equal_272_i11_2_lut_rep_73_3_lut_4_lut (.A(addr_c_2), .B(addr_c_3), 
         .C(addr_c_1), .D(addr_c_0), .Z(n15021)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam equal_272_i11_2_lut_rep_73_3_lut_4_lut.init = 16'hff7f;
    LUT4 mux_175_i1_3_lut_4_lut (.A(n15011), .B(n14997), .C(\array[84] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2729[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_175_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_175_i2_3_lut_4_lut (.A(n15011), .B(n14997), .C(\array[84] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2729[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_175_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_175_i3_3_lut_4_lut (.A(n15011), .B(n14997), .C(\array[84] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2729[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_175_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_273_i11_2_lut_rep_72_3_lut_4_lut (.A(addr_c_2), .B(addr_c_3), 
         .C(addr_c_1), .D(addr_c_0), .Z(n15020)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam equal_273_i11_2_lut_rep_72_3_lut_4_lut.init = 16'hf7ff;
    LUT4 equal_274_i11_2_lut_rep_71_3_lut_4_lut (.A(addr_c_2), .B(addr_c_3), 
         .C(addr_c_1), .D(addr_c_0), .Z(n15019)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam equal_274_i11_2_lut_rep_71_3_lut_4_lut.init = 16'hfff7;
    LUT4 mux_175_i4_3_lut_4_lut (.A(n15011), .B(n14997), .C(\array[84] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2729[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_175_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_175_i5_3_lut_4_lut (.A(n15011), .B(n14997), .C(\array[84] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2729[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_175_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4135_2_lut_rep_75_3_lut_4_lut (.A(addr_c_0), .B(addr_c_1), .C(addr_c_3), 
         .D(addr_c_2), .Z(n15023)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i4135_2_lut_rep_75_3_lut_4_lut.init = 16'h8000;
    LUT4 equal_279_i11_2_lut_rep_66_3_lut_4_lut (.A(addr_c_0), .B(addr_c_1), 
         .C(addr_c_3), .D(addr_c_2), .Z(n15014)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam equal_279_i11_2_lut_rep_66_3_lut_4_lut.init = 16'hf7ff;
    LUT4 mux_175_i6_3_lut_4_lut (.A(n15011), .B(n14997), .C(\array[84] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2729[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_175_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_175_i7_3_lut_4_lut (.A(n15011), .B(n14997), .C(\array[84] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2729[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_175_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_275_i11_2_lut_rep_70_3_lut_4_lut (.A(addr_c_0), .B(addr_c_1), 
         .C(addr_c_3), .D(addr_c_2), .Z(n15018)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam equal_275_i11_2_lut_rep_70_3_lut_4_lut.init = 16'hff7f;
    LUT4 mux_175_i8_3_lut_4_lut (.A(n15011), .B(n14997), .C(\array[84] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2729[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_175_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_174_i1_3_lut_4_lut (.A(n15012), .B(n14997), .C(\array[85] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2737[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_174_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_283_i11_2_lut_rep_62_3_lut_4_lut (.A(addr_c_0), .B(addr_c_1), 
         .C(addr_c_3), .D(addr_c_2), .Z(n15010)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam equal_283_i11_2_lut_rep_62_3_lut_4_lut.init = 16'hfff7;
    LUT4 mux_174_i2_3_lut_4_lut (.A(n15012), .B(n14997), .C(\array[85] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2737[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_174_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_174_i3_3_lut_4_lut (.A(n15012), .B(n14997), .C(\array[85] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2737[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_174_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_174_i4_3_lut_4_lut (.A(n15012), .B(n14997), .C(\array[85] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2737[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_174_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_174_i5_3_lut_4_lut (.A(n15012), .B(n14997), .C(\array[85] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2737[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_174_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_287_i14_2_lut_rep_58_3_lut_4_lut (.A(addr_c_6), .B(addr_c_7), 
         .C(addr_c_5), .D(addr_c_4), .Z(n15006)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam equal_287_i14_2_lut_rep_58_3_lut_4_lut.init = 16'hff7f;
    LUT4 mux_174_i6_3_lut_4_lut (.A(n15012), .B(n14997), .C(\array[85] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2737[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_174_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_174_i7_3_lut_4_lut (.A(n15012), .B(n14997), .C(\array[85] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2737[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_174_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_303_i14_2_lut_rep_57_3_lut_4_lut (.A(addr_c_6), .B(addr_c_7), 
         .C(addr_c_5), .D(addr_c_4), .Z(n15005)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam equal_303_i14_2_lut_rep_57_3_lut_4_lut.init = 16'hf7ff;
    LUT4 mux_174_i8_3_lut_4_lut (.A(n15012), .B(n14997), .C(\array[85] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2737[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_174_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_173_i1_3_lut_4_lut (.A(n15013), .B(n14997), .C(\array[86] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2745[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_173_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_173_i2_3_lut_4_lut (.A(n15013), .B(n14997), .C(\array[86] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2745[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_173_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_319_i14_2_lut_rep_56_3_lut_4_lut (.A(addr_c_6), .B(addr_c_7), 
         .C(addr_c_5), .D(addr_c_4), .Z(n15004)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam equal_319_i14_2_lut_rep_56_3_lut_4_lut.init = 16'hfff7;
    LUT4 equal_336_i14_2_lut_rep_55_3_lut_4_lut (.A(addr_c_4), .B(addr_c_5), 
         .C(addr_c_7), .D(addr_c_6), .Z(n15003)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam equal_336_i14_2_lut_rep_55_3_lut_4_lut.init = 16'hff7f;
    LUT4 mux_173_i3_3_lut_4_lut (.A(n15013), .B(n14997), .C(\array[86] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2745[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_173_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_173_i4_3_lut_4_lut (.A(n15013), .B(n14997), .C(\array[86] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2745[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_173_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_173_i5_3_lut_4_lut (.A(n15013), .B(n14997), .C(\array[86] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2745[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_173_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_400_i14_2_lut_rep_51_3_lut_4_lut (.A(addr_c_4), .B(addr_c_5), 
         .C(addr_c_7), .D(addr_c_6), .Z(n14999)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam equal_400_i14_2_lut_rep_51_3_lut_4_lut.init = 16'hf7ff;
    LUT4 equal_464_i14_2_lut_rep_47_3_lut_4_lut (.A(addr_c_4), .B(addr_c_5), 
         .C(addr_c_7), .D(addr_c_6), .Z(n14995)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam equal_464_i14_2_lut_rep_47_3_lut_4_lut.init = 16'hfff7;
    LUT4 mux_173_i6_3_lut_4_lut (.A(n15013), .B(n14997), .C(\array[86] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2745[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_173_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_173_i7_3_lut_4_lut (.A(n15013), .B(n14997), .C(\array[86] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2745[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_173_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4137_2_lut_rep_74_3_lut_4_lut (.A(addr_c_4), .B(addr_c_5), .C(addr_c_7), 
         .D(addr_c_6), .Z(n15022)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i4137_2_lut_rep_74_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_173_i8_3_lut_4_lut (.A(n15013), .B(n14997), .C(\array[86] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2745[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_173_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_172_i1_3_lut_4_lut (.A(n15014), .B(n14997), .C(\array[87] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2753[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_172_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_172_i2_3_lut_4_lut (.A(n15014), .B(n14997), .C(\array[87] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2753[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_172_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_172_i3_3_lut_4_lut (.A(n15014), .B(n14997), .C(\array[87] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2753[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_172_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_172_i4_3_lut_4_lut (.A(n15014), .B(n14997), .C(\array[87] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2753[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_172_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_172_i5_3_lut_4_lut (.A(n15014), .B(n14997), .C(\array[87] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2753[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_172_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_172_i6_3_lut_4_lut (.A(n15014), .B(n14997), .C(\array[87] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2753[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_172_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_172_i7_3_lut_4_lut (.A(n15014), .B(n14997), .C(\array[87] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2753[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_172_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_172_i8_3_lut_4_lut (.A(n15014), .B(n14997), .C(\array[87] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2753[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_172_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_171_i1_3_lut_4_lut (.A(n15015), .B(n14997), .C(\array[88] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2761[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_171_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_171_i2_3_lut_4_lut (.A(n15015), .B(n14997), .C(\array[88] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2761[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_171_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_171_i3_3_lut_4_lut (.A(n15015), .B(n14997), .C(\array[88] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2761[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_171_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_171_i4_3_lut_4_lut (.A(n15015), .B(n14997), .C(\array[88] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2761[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_171_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_171_i5_3_lut_4_lut (.A(n15015), .B(n14997), .C(\array[88] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2761[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_171_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_171_i6_3_lut_4_lut (.A(n15015), .B(n14997), .C(\array[88] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2761[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_171_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_171_i7_3_lut_4_lut (.A(n15015), .B(n14997), .C(\array[88] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2761[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_171_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_171_i8_3_lut_4_lut (.A(n15015), .B(n14997), .C(\array[88] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2761[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_171_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_170_i1_3_lut_4_lut (.A(n15016), .B(n14997), .C(\array[89] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2769[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_170_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_170_i2_3_lut_4_lut (.A(n15016), .B(n14997), .C(\array[89] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2769[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_170_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_170_i3_3_lut_4_lut (.A(n15016), .B(n14997), .C(\array[89] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2769[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_170_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_170_i4_3_lut_4_lut (.A(n15016), .B(n14997), .C(\array[89] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2769[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_170_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_170_i5_3_lut_4_lut (.A(n15016), .B(n14997), .C(\array[89] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2769[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_170_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_170_i6_3_lut_4_lut (.A(n15016), .B(n14997), .C(\array[89] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2769[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_170_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_170_i7_3_lut_4_lut (.A(n15016), .B(n14997), .C(\array[89] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2769[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_170_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_170_i8_3_lut_4_lut (.A(n15016), .B(n14997), .C(\array[89] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2769[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_170_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_169_i1_3_lut_4_lut (.A(n15017), .B(n14997), .C(\array[90] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2777[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_169_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_169_i2_3_lut_4_lut (.A(n15017), .B(n14997), .C(\array[90] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2777[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_169_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_169_i3_3_lut_4_lut (.A(n15017), .B(n14997), .C(\array[90] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2777[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_169_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_169_i4_3_lut_4_lut (.A(n15017), .B(n14997), .C(\array[90] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2777[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_169_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_169_i5_3_lut_4_lut (.A(n15017), .B(n14997), .C(\array[90] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2777[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_169_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_169_i6_3_lut_4_lut (.A(n15017), .B(n14997), .C(\array[90] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2777[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_169_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_169_i7_3_lut_4_lut (.A(n15017), .B(n14997), .C(\array[90] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2777[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_169_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_169_i8_3_lut_4_lut (.A(n15017), .B(n14997), .C(\array[90] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2777[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_169_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_168_i1_3_lut_4_lut (.A(n15018), .B(n14997), .C(\array[91] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2785[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_168_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_168_i2_3_lut_4_lut (.A(n15018), .B(n14997), .C(\array[91] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2785[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_168_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_168_i3_3_lut_4_lut (.A(n15018), .B(n14997), .C(\array[91] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2785[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_168_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_168_i4_3_lut_4_lut (.A(n15018), .B(n14997), .C(\array[91] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2785[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_168_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_168_i5_3_lut_4_lut (.A(n15018), .B(n14997), .C(\array[91] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2785[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_168_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_168_i6_3_lut_4_lut (.A(n15018), .B(n14997), .C(\array[91] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2785[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_168_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_168_i7_3_lut_4_lut (.A(n15018), .B(n14997), .C(\array[91] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2785[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_168_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_168_i8_3_lut_4_lut (.A(n15018), .B(n14997), .C(\array[91] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2785[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_168_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_167_i1_3_lut_4_lut (.A(n15019), .B(n14997), .C(\array[92] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2793[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_167_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_167_i2_3_lut_4_lut (.A(n15019), .B(n14997), .C(\array[92] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2793[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_167_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_167_i3_3_lut_4_lut (.A(n15019), .B(n14997), .C(\array[92] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2793[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_167_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_167_i4_3_lut_4_lut (.A(n15019), .B(n14997), .C(\array[92] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2793[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_167_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_167_i5_3_lut_4_lut (.A(n15019), .B(n14997), .C(\array[92] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2793[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_167_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_167_i6_3_lut_4_lut (.A(n15019), .B(n14997), .C(\array[92] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2793[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_167_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_167_i7_3_lut_4_lut (.A(n15019), .B(n14997), .C(\array[92] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2793[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_167_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_167_i8_3_lut_4_lut (.A(n15019), .B(n14997), .C(\array[92] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2793[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_167_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_166_i1_3_lut_4_lut (.A(n15020), .B(n14997), .C(\array[93] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2801[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_166_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_166_i2_3_lut_4_lut (.A(n15020), .B(n14997), .C(\array[93] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2801[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_166_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_166_i3_3_lut_4_lut (.A(n15020), .B(n14997), .C(\array[93] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2801[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_166_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_166_i4_3_lut_4_lut (.A(n15020), .B(n14997), .C(\array[93] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2801[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_166_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_166_i5_3_lut_4_lut (.A(n15020), .B(n14997), .C(\array[93] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2801[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_166_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_166_i6_3_lut_4_lut (.A(n15020), .B(n14997), .C(\array[93] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2801[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_166_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_166_i7_3_lut_4_lut (.A(n15020), .B(n14997), .C(\array[93] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2801[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_166_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_166_i8_3_lut_4_lut (.A(n15020), .B(n14997), .C(\array[93] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2801[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_166_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_165_i1_3_lut_4_lut (.A(n15021), .B(n14997), .C(\array[94] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2809[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_165_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_165_i2_3_lut_4_lut (.A(n15021), .B(n14997), .C(\array[94] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2809[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_165_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_165_i3_3_lut_4_lut (.A(n15021), .B(n14997), .C(\array[94] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2809[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_165_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_165_i4_3_lut_4_lut (.A(n15021), .B(n14997), .C(\array[94] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2809[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_165_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_165_i5_3_lut_4_lut (.A(n15021), .B(n14997), .C(\array[94] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2809[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_165_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_165_i6_3_lut_4_lut (.A(n15021), .B(n14997), .C(\array[94] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2809[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_165_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_165_i7_3_lut_4_lut (.A(n15021), .B(n14997), .C(\array[94] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2809[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_165_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_165_i8_3_lut_4_lut (.A(n15021), .B(n14997), .C(\array[94] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2809[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_165_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_164_i1_3_lut_4_lut (.A(n15023), .B(n14997), .C(\array[95] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2817[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_164_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_164_i2_3_lut_4_lut (.A(n15023), .B(n14997), .C(\array[95] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2817[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_164_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_164_i3_3_lut_4_lut (.A(n15023), .B(n14997), .C(\array[95] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2817[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_164_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_164_i4_3_lut_4_lut (.A(n15023), .B(n14997), .C(\array[95] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2817[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_164_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_164_i5_3_lut_4_lut (.A(n15023), .B(n14997), .C(\array[95] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2817[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_164_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_164_i6_3_lut_4_lut (.A(n15023), .B(n14997), .C(\array[95] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2817[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_164_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_164_i7_3_lut_4_lut (.A(n15023), .B(n14997), .C(\array[95] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2817[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_164_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_164_i8_3_lut_4_lut (.A(n15023), .B(n14997), .C(\array[95] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2817[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_164_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_163_i1_3_lut_4_lut (.A(n15007), .B(n14998), .C(\array[96] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2825[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_163_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_163_i2_3_lut_4_lut (.A(n15007), .B(n14998), .C(\array[96] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2825[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_163_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_163_i3_3_lut_4_lut (.A(n15007), .B(n14998), .C(\array[96] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2825[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_163_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_163_i4_3_lut_4_lut (.A(n15007), .B(n14998), .C(\array[96] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2825[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_163_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_163_i5_3_lut_4_lut (.A(n15007), .B(n14998), .C(\array[96] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2825[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_163_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_163_i6_3_lut_4_lut (.A(n15007), .B(n14998), .C(\array[96] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2825[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_163_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_163_i7_3_lut_4_lut (.A(n15007), .B(n14998), .C(\array[96] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2825[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_163_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_163_i8_3_lut_4_lut (.A(n15007), .B(n14998), .C(\array[96] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2825[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_163_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_162_i1_3_lut_4_lut (.A(n15008), .B(n14998), .C(\array[97] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2833[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_162_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_162_i2_3_lut_4_lut (.A(n15008), .B(n14998), .C(\array[97] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2833[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_162_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_162_i3_3_lut_4_lut (.A(n15008), .B(n14998), .C(\array[97] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2833[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_162_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_162_i4_3_lut_4_lut (.A(n15008), .B(n14998), .C(\array[97] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2833[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_162_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_162_i5_3_lut_4_lut (.A(n15008), .B(n14998), .C(\array[97] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2833[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_162_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_162_i6_3_lut_4_lut (.A(n15008), .B(n14998), .C(\array[97] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2833[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_162_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_162_i7_3_lut_4_lut (.A(n15008), .B(n14998), .C(\array[97] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2833[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_162_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_162_i8_3_lut_4_lut (.A(n15008), .B(n14998), .C(\array[97] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2833[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_162_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_161_i1_3_lut_4_lut (.A(n15009), .B(n14998), .C(\array[98] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2841[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_161_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_161_i2_3_lut_4_lut (.A(n15009), .B(n14998), .C(\array[98] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2841[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_161_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_161_i3_3_lut_4_lut (.A(n15009), .B(n14998), .C(\array[98] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2841[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_161_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_161_i4_3_lut_4_lut (.A(n15009), .B(n14998), .C(\array[98] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2841[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_161_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_161_i5_3_lut_4_lut (.A(n15009), .B(n14998), .C(\array[98] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2841[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_161_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_161_i6_3_lut_4_lut (.A(n15009), .B(n14998), .C(\array[98] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2841[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_161_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_161_i7_3_lut_4_lut (.A(n15009), .B(n14998), .C(\array[98] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2841[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_161_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_161_i8_3_lut_4_lut (.A(n15009), .B(n14998), .C(\array[98] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2841[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_161_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_160_i1_3_lut_4_lut (.A(n15010), .B(n14998), .C(\array[99] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2849[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_160_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_160_i2_3_lut_4_lut (.A(n15010), .B(n14998), .C(\array[99] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2849[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_160_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_160_i3_3_lut_4_lut (.A(n15010), .B(n14998), .C(\array[99] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2849[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_160_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_160_i4_3_lut_4_lut (.A(n15010), .B(n14998), .C(\array[99] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2849[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_160_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_160_i5_3_lut_4_lut (.A(n15010), .B(n14998), .C(\array[99] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2849[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_160_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_160_i6_3_lut_4_lut (.A(n15010), .B(n14998), .C(\array[99] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2849[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_160_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_160_i7_3_lut_4_lut (.A(n15010), .B(n14998), .C(\array[99] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2849[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_160_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_160_i8_3_lut_4_lut (.A(n15010), .B(n14998), .C(\array[99] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2849[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_160_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_159_i1_3_lut_4_lut (.A(n15011), .B(n14998), .C(\array[100] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2857[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_159_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_159_i2_3_lut_4_lut (.A(n15011), .B(n14998), .C(\array[100] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2857[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_159_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_159_i3_3_lut_4_lut (.A(n15011), .B(n14998), .C(\array[100] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2857[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_159_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_159_i4_3_lut_4_lut (.A(n15011), .B(n14998), .C(\array[100] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2857[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_159_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_159_i5_3_lut_4_lut (.A(n15011), .B(n14998), .C(\array[100] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2857[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_159_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_159_i6_3_lut_4_lut (.A(n15011), .B(n14998), .C(\array[100] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2857[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_159_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_159_i7_3_lut_4_lut (.A(n15011), .B(n14998), .C(\array[100] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2857[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_159_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_159_i8_3_lut_4_lut (.A(n15011), .B(n14998), .C(\array[100] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2857[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_159_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i1_3_lut_4_lut (.A(n15012), .B(n14998), .C(\array[101] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2865[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_158_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i2_3_lut_4_lut (.A(n15012), .B(n14998), .C(\array[101] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2865[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_158_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i3_3_lut_4_lut (.A(n15012), .B(n14998), .C(\array[101] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2865[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_158_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i4_3_lut_4_lut (.A(n15012), .B(n14998), .C(\array[101] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2865[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_158_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i5_3_lut_4_lut (.A(n15012), .B(n14998), .C(\array[101] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2865[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_158_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i6_3_lut_4_lut (.A(n15012), .B(n14998), .C(\array[101] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2865[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_158_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i7_3_lut_4_lut (.A(n15012), .B(n14998), .C(\array[101] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2865[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_158_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i8_3_lut_4_lut (.A(n15012), .B(n14998), .C(\array[101] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2865[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_158_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_157_i1_3_lut_4_lut (.A(n15013), .B(n14998), .C(\array[102] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2873[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_157_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_157_i2_3_lut_4_lut (.A(n15013), .B(n14998), .C(\array[102] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2873[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_157_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_157_i3_3_lut_4_lut (.A(n15013), .B(n14998), .C(\array[102] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2873[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_157_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_157_i4_3_lut_4_lut (.A(n15013), .B(n14998), .C(\array[102] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2873[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_157_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_157_i5_3_lut_4_lut (.A(n15013), .B(n14998), .C(\array[102] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2873[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_157_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_157_i6_3_lut_4_lut (.A(n15013), .B(n14998), .C(\array[102] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2873[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_157_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_157_i7_3_lut_4_lut (.A(n15013), .B(n14998), .C(\array[102] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2873[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_157_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_157_i8_3_lut_4_lut (.A(n15013), .B(n14998), .C(\array[102] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2873[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_157_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_156_i1_3_lut_4_lut (.A(n15014), .B(n14998), .C(\array[103] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2881[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_156_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_156_i2_3_lut_4_lut (.A(n15014), .B(n14998), .C(\array[103] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2881[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_156_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_156_i3_3_lut_4_lut (.A(n15014), .B(n14998), .C(\array[103] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2881[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_156_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_156_i4_3_lut_4_lut (.A(n15014), .B(n14998), .C(\array[103] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2881[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_156_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_156_i5_3_lut_4_lut (.A(n15014), .B(n14998), .C(\array[103] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2881[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_156_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_156_i6_3_lut_4_lut (.A(n15014), .B(n14998), .C(\array[103] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2881[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_156_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_156_i7_3_lut_4_lut (.A(n15014), .B(n14998), .C(\array[103] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2881[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_156_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_156_i8_3_lut_4_lut (.A(n15014), .B(n14998), .C(\array[103] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2881[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_156_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_155_i1_3_lut_4_lut (.A(n15015), .B(n14998), .C(\array[104] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2889[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_155_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_155_i2_3_lut_4_lut (.A(n15015), .B(n14998), .C(\array[104] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2889[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_155_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_155_i3_3_lut_4_lut (.A(n15015), .B(n14998), .C(\array[104] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2889[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_155_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_155_i4_3_lut_4_lut (.A(n15015), .B(n14998), .C(\array[104] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2889[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_155_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_155_i5_3_lut_4_lut (.A(n15015), .B(n14998), .C(\array[104] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2889[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_155_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_155_i6_3_lut_4_lut (.A(n15015), .B(n14998), .C(\array[104] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2889[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_155_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_155_i7_3_lut_4_lut (.A(n15015), .B(n14998), .C(\array[104] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2889[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_155_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_155_i8_3_lut_4_lut (.A(n15015), .B(n14998), .C(\array[104] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2889[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_155_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_154_i1_3_lut_4_lut (.A(n15016), .B(n14998), .C(\array[105] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2897[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_154_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_154_i2_3_lut_4_lut (.A(n15016), .B(n14998), .C(\array[105] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2897[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_154_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_154_i3_3_lut_4_lut (.A(n15016), .B(n14998), .C(\array[105] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2897[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_154_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_154_i4_3_lut_4_lut (.A(n15016), .B(n14998), .C(\array[105] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2897[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_154_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_154_i5_3_lut_4_lut (.A(n15016), .B(n14998), .C(\array[105] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2897[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_154_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_154_i6_3_lut_4_lut (.A(n15016), .B(n14998), .C(\array[105] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2897[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_154_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_154_i7_3_lut_4_lut (.A(n15016), .B(n14998), .C(\array[105] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2897[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_154_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_154_i8_3_lut_4_lut (.A(n15016), .B(n14998), .C(\array[105] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2897[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_154_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_153_i1_3_lut_4_lut (.A(n15017), .B(n14998), .C(\array[106] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2905[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_153_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_153_i2_3_lut_4_lut (.A(n15017), .B(n14998), .C(\array[106] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2905[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_153_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_153_i3_3_lut_4_lut (.A(n15017), .B(n14998), .C(\array[106] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2905[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_153_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_153_i4_3_lut_4_lut (.A(n15017), .B(n14998), .C(\array[106] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2905[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_153_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_153_i5_3_lut_4_lut (.A(n15017), .B(n14998), .C(\array[106] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2905[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_153_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_153_i6_3_lut_4_lut (.A(n15017), .B(n14998), .C(\array[106] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2905[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_153_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_153_i7_3_lut_4_lut (.A(n15017), .B(n14998), .C(\array[106] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2905[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_153_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_153_i8_3_lut_4_lut (.A(n15017), .B(n14998), .C(\array[106] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2905[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_153_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_152_i1_3_lut_4_lut (.A(n15018), .B(n14998), .C(\array[107] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2913[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_152_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_152_i2_3_lut_4_lut (.A(n15018), .B(n14998), .C(\array[107] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2913[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_152_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_152_i3_3_lut_4_lut (.A(n15018), .B(n14998), .C(\array[107] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2913[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_152_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_152_i4_3_lut_4_lut (.A(n15018), .B(n14998), .C(\array[107] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2913[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_152_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_152_i5_3_lut_4_lut (.A(n15018), .B(n14998), .C(\array[107] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2913[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_152_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_152_i6_3_lut_4_lut (.A(n15018), .B(n14998), .C(\array[107] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2913[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_152_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_152_i7_3_lut_4_lut (.A(n15018), .B(n14998), .C(\array[107] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2913[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_152_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_152_i8_3_lut_4_lut (.A(n15018), .B(n14998), .C(\array[107] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2913[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_152_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_151_i1_3_lut_4_lut (.A(n15019), .B(n14998), .C(\array[108] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2921[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_151_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_151_i2_3_lut_4_lut (.A(n15019), .B(n14998), .C(\array[108] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2921[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_151_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_151_i3_3_lut_4_lut (.A(n15019), .B(n14998), .C(\array[108] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2921[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_151_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_151_i4_3_lut_4_lut (.A(n15019), .B(n14998), .C(\array[108] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2921[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_151_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_151_i5_3_lut_4_lut (.A(n15019), .B(n14998), .C(\array[108] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2921[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_151_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_151_i6_3_lut_4_lut (.A(n15019), .B(n14998), .C(\array[108] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2921[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_151_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_151_i7_3_lut_4_lut (.A(n15019), .B(n14998), .C(\array[108] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2921[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_151_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_151_i8_3_lut_4_lut (.A(n15019), .B(n14998), .C(\array[108] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2921[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_151_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_150_i1_3_lut_4_lut (.A(n15020), .B(n14998), .C(\array[109] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2929[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_150_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_150_i2_3_lut_4_lut (.A(n15020), .B(n14998), .C(\array[109] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2929[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_150_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_150_i3_3_lut_4_lut (.A(n15020), .B(n14998), .C(\array[109] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2929[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_150_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_150_i4_3_lut_4_lut (.A(n15020), .B(n14998), .C(\array[109] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2929[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_150_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_150_i5_3_lut_4_lut (.A(n15020), .B(n14998), .C(\array[109] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2929[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_150_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_150_i6_3_lut_4_lut (.A(n15020), .B(n14998), .C(\array[109] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2929[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_150_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_150_i7_3_lut_4_lut (.A(n15020), .B(n14998), .C(\array[109] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2929[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_150_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_150_i8_3_lut_4_lut (.A(n15020), .B(n14998), .C(\array[109] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2929[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_150_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_149_i1_3_lut_4_lut (.A(n15021), .B(n14998), .C(\array[110] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2937[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_149_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_149_i2_3_lut_4_lut (.A(n15021), .B(n14998), .C(\array[110] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2937[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_149_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_149_i3_3_lut_4_lut (.A(n15021), .B(n14998), .C(\array[110] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2937[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_149_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_149_i4_3_lut_4_lut (.A(n15021), .B(n14998), .C(\array[110] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2937[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_149_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_149_i5_3_lut_4_lut (.A(n15021), .B(n14998), .C(\array[110] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2937[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_149_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_149_i6_3_lut_4_lut (.A(n15021), .B(n14998), .C(\array[110] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2937[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_149_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_149_i7_3_lut_4_lut (.A(n15021), .B(n14998), .C(\array[110] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2937[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_149_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_149_i8_3_lut_4_lut (.A(n15021), .B(n14998), .C(\array[110] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2937[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_149_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_148_i1_3_lut_4_lut (.A(n15023), .B(n14998), .C(\array[111] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2945[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_148_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_148_i2_3_lut_4_lut (.A(n15023), .B(n14998), .C(\array[111] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2945[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_148_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_148_i3_3_lut_4_lut (.A(n15023), .B(n14998), .C(\array[111] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2945[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_148_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_148_i4_3_lut_4_lut (.A(n15023), .B(n14998), .C(\array[111] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2945[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_148_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_148_i5_3_lut_4_lut (.A(n15023), .B(n14998), .C(\array[111] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2945[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_148_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_148_i6_3_lut_4_lut (.A(n15023), .B(n14998), .C(\array[111] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2945[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_148_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_148_i7_3_lut_4_lut (.A(n15023), .B(n14998), .C(\array[111] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2945[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_148_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_148_i8_3_lut_4_lut (.A(n15023), .B(n14998), .C(\array[111] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2945[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_148_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_147_i1_3_lut_4_lut (.A(n15007), .B(n14999), .C(\array[112] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2953[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_147_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_147_i2_3_lut_4_lut (.A(n15007), .B(n14999), .C(\array[112] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2953[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_147_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_147_i3_3_lut_4_lut (.A(n15007), .B(n14999), .C(\array[112] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2953[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_147_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_147_i4_3_lut_4_lut (.A(n15007), .B(n14999), .C(\array[112] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2953[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_147_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_147_i5_3_lut_4_lut (.A(n15007), .B(n14999), .C(\array[112] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2953[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_147_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_147_i6_3_lut_4_lut (.A(n15007), .B(n14999), .C(\array[112] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2953[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_147_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_147_i7_3_lut_4_lut (.A(n15007), .B(n14999), .C(\array[112] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2953[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_147_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_147_i8_3_lut_4_lut (.A(n15007), .B(n14999), .C(\array[112] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2953[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_147_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_146_i1_3_lut_4_lut (.A(n15008), .B(n14999), .C(\array[113] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2961[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_146_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_146_i2_3_lut_4_lut (.A(n15008), .B(n14999), .C(\array[113] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2961[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_146_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_146_i3_3_lut_4_lut (.A(n15008), .B(n14999), .C(\array[113] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2961[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_146_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_146_i4_3_lut_4_lut (.A(n15008), .B(n14999), .C(\array[113] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2961[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_146_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_146_i5_3_lut_4_lut (.A(n15008), .B(n14999), .C(\array[113] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2961[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_146_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_146_i6_3_lut_4_lut (.A(n15008), .B(n14999), .C(\array[113] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2961[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_146_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_146_i7_3_lut_4_lut (.A(n15008), .B(n14999), .C(\array[113] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2961[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_146_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_146_i8_3_lut_4_lut (.A(n15008), .B(n14999), .C(\array[113] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2961[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_146_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_145_i1_3_lut_4_lut (.A(n15009), .B(n14999), .C(\array[114] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2969[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_145_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_145_i2_3_lut_4_lut (.A(n15009), .B(n14999), .C(\array[114] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2969[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_145_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_145_i3_3_lut_4_lut (.A(n15009), .B(n14999), .C(\array[114] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2969[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_145_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_145_i4_3_lut_4_lut (.A(n15009), .B(n14999), .C(\array[114] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2969[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_145_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_145_i5_3_lut_4_lut (.A(n15009), .B(n14999), .C(\array[114] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2969[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_145_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_145_i6_3_lut_4_lut (.A(n15009), .B(n14999), .C(\array[114] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2969[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_145_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_145_i7_3_lut_4_lut (.A(n15009), .B(n14999), .C(\array[114] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2969[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_145_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_145_i8_3_lut_4_lut (.A(n15009), .B(n14999), .C(\array[114] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2969[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_145_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_144_i1_3_lut_4_lut (.A(n15010), .B(n14999), .C(\array[115] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2977[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_144_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_144_i2_3_lut_4_lut (.A(n15010), .B(n14999), .C(\array[115] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2977[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_144_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_144_i3_3_lut_4_lut (.A(n15010), .B(n14999), .C(\array[115] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2977[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_144_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_144_i4_3_lut_4_lut (.A(n15010), .B(n14999), .C(\array[115] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2977[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_144_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_144_i5_3_lut_4_lut (.A(n15010), .B(n14999), .C(\array[115] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2977[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_144_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_144_i6_3_lut_4_lut (.A(n15010), .B(n14999), .C(\array[115] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2977[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_144_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_144_i7_3_lut_4_lut (.A(n15010), .B(n14999), .C(\array[115] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2977[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_144_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_144_i8_3_lut_4_lut (.A(n15010), .B(n14999), .C(\array[115] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2977[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_144_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_143_i1_3_lut_4_lut (.A(n15011), .B(n14999), .C(\array[116] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2985[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_143_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_143_i2_3_lut_4_lut (.A(n15011), .B(n14999), .C(\array[116] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2985[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_143_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_143_i3_3_lut_4_lut (.A(n15011), .B(n14999), .C(\array[116] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2985[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_143_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_143_i4_3_lut_4_lut (.A(n15011), .B(n14999), .C(\array[116] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2985[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_143_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_143_i5_3_lut_4_lut (.A(n15011), .B(n14999), .C(\array[116] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2985[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_143_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_143_i6_3_lut_4_lut (.A(n15011), .B(n14999), .C(\array[116] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2985[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_143_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_143_i7_3_lut_4_lut (.A(n15011), .B(n14999), .C(\array[116] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2985[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_143_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_143_i8_3_lut_4_lut (.A(n15011), .B(n14999), .C(\array[116] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2985[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_143_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_142_i1_3_lut_4_lut (.A(n15012), .B(n14999), .C(\array[117] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2993[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_142_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_142_i2_3_lut_4_lut (.A(n15012), .B(n14999), .C(\array[117] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2993[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_142_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_142_i3_3_lut_4_lut (.A(n15012), .B(n14999), .C(\array[117] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2993[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_142_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_142_i4_3_lut_4_lut (.A(n15012), .B(n14999), .C(\array[117] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2993[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_142_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_142_i5_3_lut_4_lut (.A(n15012), .B(n14999), .C(\array[117] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2993[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_142_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_142_i6_3_lut_4_lut (.A(n15012), .B(n14999), .C(\array[117] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2993[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_142_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_142_i7_3_lut_4_lut (.A(n15012), .B(n14999), .C(\array[117] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2993[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_142_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_142_i8_3_lut_4_lut (.A(n15012), .B(n14999), .C(\array[117] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2993[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_142_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_141_i1_3_lut_4_lut (.A(n15013), .B(n14999), .C(\array[118] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3001[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_141_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_141_i2_3_lut_4_lut (.A(n15013), .B(n14999), .C(\array[118] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3001[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_141_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_141_i3_3_lut_4_lut (.A(n15013), .B(n14999), .C(\array[118] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3001[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_141_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_255_i4_3_lut_4_lut (.A(n15011), .B(n14992), .C(\array[4] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2089[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_255_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_141_i4_3_lut_4_lut (.A(n15013), .B(n14999), .C(\array[118] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3001[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_141_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_141_i5_3_lut_4_lut (.A(n15013), .B(n14999), .C(\array[118] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3001[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_141_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_141_i6_3_lut_4_lut (.A(n15013), .B(n14999), .C(\array[118] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3001[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_141_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_141_i7_3_lut_4_lut (.A(n15013), .B(n14999), .C(\array[118] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3001[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_141_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_141_i8_3_lut_4_lut (.A(n15013), .B(n14999), .C(\array[118] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3001[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_141_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_140_i1_3_lut_4_lut (.A(n15014), .B(n14999), .C(\array[119] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3009[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_140_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_140_i2_3_lut_4_lut (.A(n15014), .B(n14999), .C(\array[119] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3009[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_140_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_140_i3_3_lut_4_lut (.A(n15014), .B(n14999), .C(\array[119] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3009[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_140_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_140_i4_3_lut_4_lut (.A(n15014), .B(n14999), .C(\array[119] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3009[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_140_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_140_i5_3_lut_4_lut (.A(n15014), .B(n14999), .C(\array[119] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3009[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_140_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_140_i6_3_lut_4_lut (.A(n15014), .B(n14999), .C(\array[119] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3009[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_140_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_140_i7_3_lut_4_lut (.A(n15014), .B(n14999), .C(\array[119] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3009[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_140_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_140_i8_3_lut_4_lut (.A(n15014), .B(n14999), .C(\array[119] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3009[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_140_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_139_i1_3_lut_4_lut (.A(n15015), .B(n14999), .C(\array[120] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3017[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_139_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_139_i2_3_lut_4_lut (.A(n15015), .B(n14999), .C(\array[120] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3017[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_139_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_139_i3_3_lut_4_lut (.A(n15015), .B(n14999), .C(\array[120] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3017[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_139_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_139_i4_3_lut_4_lut (.A(n15015), .B(n14999), .C(\array[120] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3017[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_139_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_139_i5_3_lut_4_lut (.A(n15015), .B(n14999), .C(\array[120] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3017[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_139_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_139_i6_3_lut_4_lut (.A(n15015), .B(n14999), .C(\array[120] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3017[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_139_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_139_i7_3_lut_4_lut (.A(n15015), .B(n14999), .C(\array[120] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3017[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_139_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_139_i8_3_lut_4_lut (.A(n15015), .B(n14999), .C(\array[120] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3017[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_139_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_138_i1_3_lut_4_lut (.A(n15016), .B(n14999), .C(\array[121] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3025[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_138_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_138_i2_3_lut_4_lut (.A(n15016), .B(n14999), .C(\array[121] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3025[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_138_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_138_i3_3_lut_4_lut (.A(n15016), .B(n14999), .C(\array[121] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3025[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_138_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_138_i4_3_lut_4_lut (.A(n15016), .B(n14999), .C(\array[121] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3025[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_138_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_138_i5_3_lut_4_lut (.A(n15016), .B(n14999), .C(\array[121] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3025[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_138_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_138_i6_3_lut_4_lut (.A(n15016), .B(n14999), .C(\array[121] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3025[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_138_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_138_i7_3_lut_4_lut (.A(n15016), .B(n14999), .C(\array[121] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3025[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_138_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_138_i8_3_lut_4_lut (.A(n15016), .B(n14999), .C(\array[121] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3025[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_138_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_137_i1_3_lut_4_lut (.A(n15017), .B(n14999), .C(\array[122] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3033[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_137_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_137_i2_3_lut_4_lut (.A(n15017), .B(n14999), .C(\array[122] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3033[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_137_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_137_i3_3_lut_4_lut (.A(n15017), .B(n14999), .C(\array[122] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3033[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_137_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_137_i4_3_lut_4_lut (.A(n15017), .B(n14999), .C(\array[122] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3033[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_137_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_137_i5_3_lut_4_lut (.A(n15017), .B(n14999), .C(\array[122] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3033[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_137_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_137_i6_3_lut_4_lut (.A(n15017), .B(n14999), .C(\array[122] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3033[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_137_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_137_i7_3_lut_4_lut (.A(n15017), .B(n14999), .C(\array[122] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3033[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_137_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_137_i8_3_lut_4_lut (.A(n15017), .B(n14999), .C(\array[122] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3033[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_137_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_136_i1_3_lut_4_lut (.A(n15018), .B(n14999), .C(\array[123] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3041[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_136_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_136_i2_3_lut_4_lut (.A(n15018), .B(n14999), .C(\array[123] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3041[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_136_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_136_i3_3_lut_4_lut (.A(n15018), .B(n14999), .C(\array[123] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3041[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_136_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_136_i4_3_lut_4_lut (.A(n15018), .B(n14999), .C(\array[123] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3041[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_136_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_136_i5_3_lut_4_lut (.A(n15018), .B(n14999), .C(\array[123] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3041[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_136_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_136_i6_3_lut_4_lut (.A(n15018), .B(n14999), .C(\array[123] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3041[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_136_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_136_i7_3_lut_4_lut (.A(n15018), .B(n14999), .C(\array[123] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3041[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_136_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_136_i8_3_lut_4_lut (.A(n15018), .B(n14999), .C(\array[123] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3041[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_136_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_135_i1_3_lut_4_lut (.A(n15019), .B(n14999), .C(\array[124] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3049[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_135_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_135_i2_3_lut_4_lut (.A(n15019), .B(n14999), .C(\array[124] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3049[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_135_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_135_i3_3_lut_4_lut (.A(n15019), .B(n14999), .C(\array[124] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3049[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_135_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_135_i4_3_lut_4_lut (.A(n15019), .B(n14999), .C(\array[124] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3049[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_135_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_135_i5_3_lut_4_lut (.A(n15019), .B(n14999), .C(\array[124] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3049[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_135_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_135_i6_3_lut_4_lut (.A(n15019), .B(n14999), .C(\array[124] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3049[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_135_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_135_i7_3_lut_4_lut (.A(n15019), .B(n14999), .C(\array[124] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3049[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_135_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_135_i8_3_lut_4_lut (.A(n15019), .B(n14999), .C(\array[124] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3049[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_135_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_134_i1_3_lut_4_lut (.A(n15020), .B(n14999), .C(\array[125] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3057[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_134_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_134_i2_3_lut_4_lut (.A(n15020), .B(n14999), .C(\array[125] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3057[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_134_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_134_i3_3_lut_4_lut (.A(n15020), .B(n14999), .C(\array[125] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3057[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_134_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_134_i4_3_lut_4_lut (.A(n15020), .B(n14999), .C(\array[125] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3057[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_134_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_134_i5_3_lut_4_lut (.A(n15020), .B(n14999), .C(\array[125] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3057[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_134_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_134_i6_3_lut_4_lut (.A(n15020), .B(n14999), .C(\array[125] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3057[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_134_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_134_i7_3_lut_4_lut (.A(n15020), .B(n14999), .C(\array[125] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3057[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_134_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_134_i8_3_lut_4_lut (.A(n15020), .B(n14999), .C(\array[125] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3057[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_134_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_133_i1_3_lut_4_lut (.A(n15021), .B(n14999), .C(\array[126] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3065[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_133_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_133_i2_3_lut_4_lut (.A(n15021), .B(n14999), .C(\array[126] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3065[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_133_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_133_i3_3_lut_4_lut (.A(n15021), .B(n14999), .C(\array[126] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3065[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_133_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_133_i4_3_lut_4_lut (.A(n15021), .B(n14999), .C(\array[126] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3065[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_133_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_133_i5_3_lut_4_lut (.A(n15021), .B(n14999), .C(\array[126] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3065[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_133_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_133_i6_3_lut_4_lut (.A(n15021), .B(n14999), .C(\array[126] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3065[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_133_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_133_i7_3_lut_4_lut (.A(n15021), .B(n14999), .C(\array[126] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3065[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_133_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_133_i8_3_lut_4_lut (.A(n15021), .B(n14999), .C(\array[126] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3065[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_133_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_132_i1_3_lut_4_lut (.A(n15023), .B(n14999), .C(\array[127] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3073[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_132_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_132_i2_3_lut_4_lut (.A(n15023), .B(n14999), .C(\array[127] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3073[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_132_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_132_i3_3_lut_4_lut (.A(n15023), .B(n14999), .C(\array[127] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3073[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_132_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_132_i4_3_lut_4_lut (.A(n15023), .B(n14999), .C(\array[127] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3073[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_132_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_132_i5_3_lut_4_lut (.A(n15023), .B(n14999), .C(\array[127] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3073[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_132_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_132_i6_3_lut_4_lut (.A(n15023), .B(n14999), .C(\array[127] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3073[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_132_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_132_i7_3_lut_4_lut (.A(n15023), .B(n14999), .C(\array[127] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3073[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_132_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_132_i8_3_lut_4_lut (.A(n15023), .B(n14999), .C(\array[127] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3073[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_132_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_131_i1_3_lut_4_lut (.A(n15007), .B(n15000), .C(\array[128] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3081[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_131_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_131_i2_3_lut_4_lut (.A(n15007), .B(n15000), .C(\array[128] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3081[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_131_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_131_i3_3_lut_4_lut (.A(n15007), .B(n15000), .C(\array[128] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3081[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_131_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_131_i4_3_lut_4_lut (.A(n15007), .B(n15000), .C(\array[128] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3081[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_131_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_131_i5_3_lut_4_lut (.A(n15007), .B(n15000), .C(\array[128] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3081[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_131_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_131_i6_3_lut_4_lut (.A(n15007), .B(n15000), .C(\array[128] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3081[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_131_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_131_i7_3_lut_4_lut (.A(n15007), .B(n15000), .C(\array[128] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3081[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_131_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_131_i8_3_lut_4_lut (.A(n15007), .B(n15000), .C(\array[128] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3081[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_131_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_130_i1_3_lut_4_lut (.A(n15008), .B(n15000), .C(\array[129] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3089[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_130_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_130_i2_3_lut_4_lut (.A(n15008), .B(n15000), .C(\array[129] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3089[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_130_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_130_i3_3_lut_4_lut (.A(n15008), .B(n15000), .C(\array[129] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3089[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_130_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_130_i4_3_lut_4_lut (.A(n15008), .B(n15000), .C(\array[129] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3089[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_130_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_130_i5_3_lut_4_lut (.A(n15008), .B(n15000), .C(\array[129] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3089[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_130_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_130_i6_3_lut_4_lut (.A(n15008), .B(n15000), .C(\array[129] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3089[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_130_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_130_i7_3_lut_4_lut (.A(n15008), .B(n15000), .C(\array[129] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3089[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_130_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_130_i8_3_lut_4_lut (.A(n15008), .B(n15000), .C(\array[129] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3089[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_130_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_129_i1_3_lut_4_lut (.A(n15009), .B(n15000), .C(\array[130] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3097[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_129_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_129_i2_3_lut_4_lut (.A(n15009), .B(n15000), .C(\array[130] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3097[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_129_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_129_i3_3_lut_4_lut (.A(n15009), .B(n15000), .C(\array[130] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3097[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_129_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_129_i4_3_lut_4_lut (.A(n15009), .B(n15000), .C(\array[130] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3097[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_129_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_129_i5_3_lut_4_lut (.A(n15009), .B(n15000), .C(\array[130] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3097[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_129_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_129_i6_3_lut_4_lut (.A(n15009), .B(n15000), .C(\array[130] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3097[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_129_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_129_i7_3_lut_4_lut (.A(n15009), .B(n15000), .C(\array[130] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3097[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_129_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_129_i8_3_lut_4_lut (.A(n15009), .B(n15000), .C(\array[130] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3097[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_129_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_128_i1_3_lut_4_lut (.A(n15010), .B(n15000), .C(\array[131] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3105[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_128_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_128_i2_3_lut_4_lut (.A(n15010), .B(n15000), .C(\array[131] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3105[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_128_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_128_i3_3_lut_4_lut (.A(n15010), .B(n15000), .C(\array[131] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3105[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_128_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_128_i4_3_lut_4_lut (.A(n15010), .B(n15000), .C(\array[131] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3105[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_128_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_128_i5_3_lut_4_lut (.A(n15010), .B(n15000), .C(\array[131] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3105[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_128_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_128_i6_3_lut_4_lut (.A(n15010), .B(n15000), .C(\array[131] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3105[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_128_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_128_i7_3_lut_4_lut (.A(n15010), .B(n15000), .C(\array[131] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3105[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_128_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_128_i8_3_lut_4_lut (.A(n15010), .B(n15000), .C(\array[131] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3105[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_128_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_127_i1_3_lut_4_lut (.A(n15011), .B(n15000), .C(\array[132] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3113[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_127_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_127_i2_3_lut_4_lut (.A(n15011), .B(n15000), .C(\array[132] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3113[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_127_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_127_i3_3_lut_4_lut (.A(n15011), .B(n15000), .C(\array[132] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3113[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_127_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_127_i4_3_lut_4_lut (.A(n15011), .B(n15000), .C(\array[132] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3113[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_127_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_127_i5_3_lut_4_lut (.A(n15011), .B(n15000), .C(\array[132] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3113[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_127_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_127_i6_3_lut_4_lut (.A(n15011), .B(n15000), .C(\array[132] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3113[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_127_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_127_i7_3_lut_4_lut (.A(n15011), .B(n15000), .C(\array[132] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3113[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_127_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_127_i8_3_lut_4_lut (.A(n15011), .B(n15000), .C(\array[132] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3113[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_127_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_126_i1_3_lut_4_lut (.A(n15012), .B(n15000), .C(\array[133] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3121[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_126_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_126_i2_3_lut_4_lut (.A(n15012), .B(n15000), .C(\array[133] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3121[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_126_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_126_i3_3_lut_4_lut (.A(n15012), .B(n15000), .C(\array[133] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3121[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_126_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_126_i4_3_lut_4_lut (.A(n15012), .B(n15000), .C(\array[133] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3121[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_126_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_126_i5_3_lut_4_lut (.A(n15012), .B(n15000), .C(\array[133] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3121[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_126_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_126_i6_3_lut_4_lut (.A(n15012), .B(n15000), .C(\array[133] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3121[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_126_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_126_i7_3_lut_4_lut (.A(n15012), .B(n15000), .C(\array[133] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3121[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_126_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_126_i8_3_lut_4_lut (.A(n15012), .B(n15000), .C(\array[133] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3121[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_126_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_125_i1_3_lut_4_lut (.A(n15013), .B(n15000), .C(\array[134] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3129[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_125_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_125_i2_3_lut_4_lut (.A(n15013), .B(n15000), .C(\array[134] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3129[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_125_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_125_i3_3_lut_4_lut (.A(n15013), .B(n15000), .C(\array[134] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3129[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_125_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_125_i4_3_lut_4_lut (.A(n15013), .B(n15000), .C(\array[134] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3129[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_125_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_125_i5_3_lut_4_lut (.A(n15013), .B(n15000), .C(\array[134] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3129[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_125_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_125_i6_3_lut_4_lut (.A(n15013), .B(n15000), .C(\array[134] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3129[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_125_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_125_i7_3_lut_4_lut (.A(n15013), .B(n15000), .C(\array[134] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3129[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_125_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_125_i8_3_lut_4_lut (.A(n15013), .B(n15000), .C(\array[134] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3129[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_125_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_124_i1_3_lut_4_lut (.A(n15014), .B(n15000), .C(\array[135] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3137[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_124_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_124_i2_3_lut_4_lut (.A(n15014), .B(n15000), .C(\array[135] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3137[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_124_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_124_i3_3_lut_4_lut (.A(n15014), .B(n15000), .C(\array[135] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3137[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_124_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_124_i4_3_lut_4_lut (.A(n15014), .B(n15000), .C(\array[135] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3137[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_124_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_124_i5_3_lut_4_lut (.A(n15014), .B(n15000), .C(\array[135] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3137[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_124_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_124_i6_3_lut_4_lut (.A(n15014), .B(n15000), .C(\array[135] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3137[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_124_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_124_i7_3_lut_4_lut (.A(n15014), .B(n15000), .C(\array[135] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3137[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_124_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_124_i8_3_lut_4_lut (.A(n15014), .B(n15000), .C(\array[135] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3137[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_124_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_123_i1_3_lut_4_lut (.A(n15015), .B(n15000), .C(\array[136] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3145[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_123_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_123_i2_3_lut_4_lut (.A(n15015), .B(n15000), .C(\array[136] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3145[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_123_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_123_i3_3_lut_4_lut (.A(n15015), .B(n15000), .C(\array[136] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3145[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_123_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_123_i4_3_lut_4_lut (.A(n15015), .B(n15000), .C(\array[136] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3145[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_123_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_123_i5_3_lut_4_lut (.A(n15015), .B(n15000), .C(\array[136] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3145[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_123_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_123_i6_3_lut_4_lut (.A(n15015), .B(n15000), .C(\array[136] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3145[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_123_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_123_i7_3_lut_4_lut (.A(n15015), .B(n15000), .C(\array[136] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3145[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_123_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_123_i8_3_lut_4_lut (.A(n15015), .B(n15000), .C(\array[136] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3145[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_123_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_122_i1_3_lut_4_lut (.A(n15016), .B(n15000), .C(\array[137] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3153[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_122_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_122_i2_3_lut_4_lut (.A(n15016), .B(n15000), .C(\array[137] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3153[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_122_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_122_i3_3_lut_4_lut (.A(n15016), .B(n15000), .C(\array[137] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3153[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_122_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_122_i4_3_lut_4_lut (.A(n15016), .B(n15000), .C(\array[137] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3153[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_122_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_122_i5_3_lut_4_lut (.A(n15016), .B(n15000), .C(\array[137] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3153[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_122_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_122_i6_3_lut_4_lut (.A(n15016), .B(n15000), .C(\array[137] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3153[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_122_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_122_i7_3_lut_4_lut (.A(n15016), .B(n15000), .C(\array[137] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3153[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_122_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_122_i8_3_lut_4_lut (.A(n15016), .B(n15000), .C(\array[137] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3153[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_122_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_121_i1_3_lut_4_lut (.A(n15017), .B(n15000), .C(\array[138] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3161[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_121_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_121_i2_3_lut_4_lut (.A(n15017), .B(n15000), .C(\array[138] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3161[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_121_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_121_i3_3_lut_4_lut (.A(n15017), .B(n15000), .C(\array[138] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3161[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_121_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_121_i4_3_lut_4_lut (.A(n15017), .B(n15000), .C(\array[138] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3161[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_121_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_121_i5_3_lut_4_lut (.A(n15017), .B(n15000), .C(\array[138] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3161[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_121_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_121_i6_3_lut_4_lut (.A(n15017), .B(n15000), .C(\array[138] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3161[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_121_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_121_i7_3_lut_4_lut (.A(n15017), .B(n15000), .C(\array[138] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3161[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_121_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_121_i8_3_lut_4_lut (.A(n15017), .B(n15000), .C(\array[138] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3161[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_121_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_120_i1_3_lut_4_lut (.A(n15018), .B(n15000), .C(\array[139] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3169[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_120_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_120_i2_3_lut_4_lut (.A(n15018), .B(n15000), .C(\array[139] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3169[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_120_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_120_i3_3_lut_4_lut (.A(n15018), .B(n15000), .C(\array[139] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3169[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_120_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_120_i4_3_lut_4_lut (.A(n15018), .B(n15000), .C(\array[139] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3169[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_120_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_120_i5_3_lut_4_lut (.A(n15018), .B(n15000), .C(\array[139] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3169[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_120_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_120_i6_3_lut_4_lut (.A(n15018), .B(n15000), .C(\array[139] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3169[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_120_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_120_i7_3_lut_4_lut (.A(n15018), .B(n15000), .C(\array[139] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3169[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_120_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_120_i8_3_lut_4_lut (.A(n15018), .B(n15000), .C(\array[139] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3169[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_120_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_119_i1_3_lut_4_lut (.A(n15019), .B(n15000), .C(\array[140] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3177[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_119_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_119_i2_3_lut_4_lut (.A(n15019), .B(n15000), .C(\array[140] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3177[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_119_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_119_i3_3_lut_4_lut (.A(n15019), .B(n15000), .C(\array[140] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3177[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_119_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_119_i4_3_lut_4_lut (.A(n15019), .B(n15000), .C(\array[140] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3177[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_119_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_119_i5_3_lut_4_lut (.A(n15019), .B(n15000), .C(\array[140] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3177[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_119_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_119_i6_3_lut_4_lut (.A(n15019), .B(n15000), .C(\array[140] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3177[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_119_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_119_i7_3_lut_4_lut (.A(n15019), .B(n15000), .C(\array[140] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3177[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_119_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_119_i8_3_lut_4_lut (.A(n15019), .B(n15000), .C(\array[140] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3177[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_119_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_118_i1_3_lut_4_lut (.A(n15020), .B(n15000), .C(\array[141] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3185[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_118_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_118_i2_3_lut_4_lut (.A(n15020), .B(n15000), .C(\array[141] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3185[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_118_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_118_i3_3_lut_4_lut (.A(n15020), .B(n15000), .C(\array[141] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3185[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_118_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_118_i4_3_lut_4_lut (.A(n15020), .B(n15000), .C(\array[141] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3185[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_118_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_118_i5_3_lut_4_lut (.A(n15020), .B(n15000), .C(\array[141] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3185[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_118_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_118_i6_3_lut_4_lut (.A(n15020), .B(n15000), .C(\array[141] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3185[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_118_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_118_i7_3_lut_4_lut (.A(n15020), .B(n15000), .C(\array[141] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3185[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_118_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_118_i8_3_lut_4_lut (.A(n15020), .B(n15000), .C(\array[141] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3185[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_118_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_117_i1_3_lut_4_lut (.A(n15021), .B(n15000), .C(\array[142] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3193[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_117_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_117_i2_3_lut_4_lut (.A(n15021), .B(n15000), .C(\array[142] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3193[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_117_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_117_i3_3_lut_4_lut (.A(n15021), .B(n15000), .C(\array[142] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3193[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_117_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_117_i4_3_lut_4_lut (.A(n15021), .B(n15000), .C(\array[142] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3193[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_117_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_117_i5_3_lut_4_lut (.A(n15021), .B(n15000), .C(\array[142] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3193[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_117_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_117_i6_3_lut_4_lut (.A(n15021), .B(n15000), .C(\array[142] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3193[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_117_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_117_i7_3_lut_4_lut (.A(n15021), .B(n15000), .C(\array[142] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3193[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_117_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_117_i8_3_lut_4_lut (.A(n15021), .B(n15000), .C(\array[142] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3193[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_117_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_116_i1_3_lut_4_lut (.A(n15023), .B(n15000), .C(\array[143] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3201[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_116_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_116_i2_3_lut_4_lut (.A(n15023), .B(n15000), .C(\array[143] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3201[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_116_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_116_i3_3_lut_4_lut (.A(n15023), .B(n15000), .C(\array[143] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3201[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_116_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_116_i4_3_lut_4_lut (.A(n15023), .B(n15000), .C(\array[143] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3201[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_116_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_116_i5_3_lut_4_lut (.A(n15023), .B(n15000), .C(\array[143] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3201[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_116_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_116_i6_3_lut_4_lut (.A(n15023), .B(n15000), .C(\array[143] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3201[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_116_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_116_i7_3_lut_4_lut (.A(n15023), .B(n15000), .C(\array[143] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3201[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_116_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_116_i8_3_lut_4_lut (.A(n15023), .B(n15000), .C(\array[143] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3201[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_116_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_115_i1_3_lut_4_lut (.A(n15007), .B(n15001), .C(\array[144] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3209[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_115_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_115_i2_3_lut_4_lut (.A(n15007), .B(n15001), .C(\array[144] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3209[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_115_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_115_i3_3_lut_4_lut (.A(n15007), .B(n15001), .C(\array[144] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3209[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_115_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_115_i4_3_lut_4_lut (.A(n15007), .B(n15001), .C(\array[144] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3209[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_115_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_115_i5_3_lut_4_lut (.A(n15007), .B(n15001), .C(\array[144] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3209[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_115_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_115_i6_3_lut_4_lut (.A(n15007), .B(n15001), .C(\array[144] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3209[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_115_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_115_i7_3_lut_4_lut (.A(n15007), .B(n15001), .C(\array[144] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3209[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_115_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_115_i8_3_lut_4_lut (.A(n15007), .B(n15001), .C(\array[144] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3209[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_115_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_114_i1_3_lut_4_lut (.A(n15008), .B(n15001), .C(\array[145] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3217[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_114_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_114_i2_3_lut_4_lut (.A(n15008), .B(n15001), .C(\array[145] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3217[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_114_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_114_i3_3_lut_4_lut (.A(n15008), .B(n15001), .C(\array[145] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3217[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_114_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_114_i4_3_lut_4_lut (.A(n15008), .B(n15001), .C(\array[145] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3217[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_114_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_114_i5_3_lut_4_lut (.A(n15008), .B(n15001), .C(\array[145] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3217[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_114_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_114_i6_3_lut_4_lut (.A(n15008), .B(n15001), .C(\array[145] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3217[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_114_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_114_i7_3_lut_4_lut (.A(n15008), .B(n15001), .C(\array[145] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3217[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_114_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_114_i8_3_lut_4_lut (.A(n15008), .B(n15001), .C(\array[145] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3217[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_114_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_113_i1_3_lut_4_lut (.A(n15009), .B(n15001), .C(\array[146] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3225[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_113_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_113_i2_3_lut_4_lut (.A(n15009), .B(n15001), .C(\array[146] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3225[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_113_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_113_i3_3_lut_4_lut (.A(n15009), .B(n15001), .C(\array[146] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3225[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_113_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_113_i4_3_lut_4_lut (.A(n15009), .B(n15001), .C(\array[146] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3225[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_113_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_113_i5_3_lut_4_lut (.A(n15009), .B(n15001), .C(\array[146] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3225[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_113_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_113_i6_3_lut_4_lut (.A(n15009), .B(n15001), .C(\array[146] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3225[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_113_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_113_i7_3_lut_4_lut (.A(n15009), .B(n15001), .C(\array[146] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3225[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_113_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_113_i8_3_lut_4_lut (.A(n15009), .B(n15001), .C(\array[146] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3225[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_113_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_112_i1_3_lut_4_lut (.A(n15010), .B(n15001), .C(\array[147] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3233[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_112_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_112_i2_3_lut_4_lut (.A(n15010), .B(n15001), .C(\array[147] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3233[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_112_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_112_i3_3_lut_4_lut (.A(n15010), .B(n15001), .C(\array[147] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3233[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_112_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_112_i4_3_lut_4_lut (.A(n15010), .B(n15001), .C(\array[147] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3233[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_112_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_112_i5_3_lut_4_lut (.A(n15010), .B(n15001), .C(\array[147] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3233[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_112_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_112_i6_3_lut_4_lut (.A(n15010), .B(n15001), .C(\array[147] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3233[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_112_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_112_i7_3_lut_4_lut (.A(n15010), .B(n15001), .C(\array[147] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3233[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_112_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_112_i8_3_lut_4_lut (.A(n15010), .B(n15001), .C(\array[147] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3233[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_112_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_111_i1_3_lut_4_lut (.A(n15011), .B(n15001), .C(\array[148] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3241[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_111_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_111_i2_3_lut_4_lut (.A(n15011), .B(n15001), .C(\array[148] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3241[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_111_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_111_i3_3_lut_4_lut (.A(n15011), .B(n15001), .C(\array[148] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3241[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_111_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_111_i4_3_lut_4_lut (.A(n15011), .B(n15001), .C(\array[148] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3241[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_111_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_111_i5_3_lut_4_lut (.A(n15011), .B(n15001), .C(\array[148] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3241[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_111_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_111_i6_3_lut_4_lut (.A(n15011), .B(n15001), .C(\array[148] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3241[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_111_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_111_i7_3_lut_4_lut (.A(n15011), .B(n15001), .C(\array[148] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3241[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_111_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_111_i8_3_lut_4_lut (.A(n15011), .B(n15001), .C(\array[148] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3241[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_111_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_110_i1_3_lut_4_lut (.A(n15012), .B(n15001), .C(\array[149] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3249[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_110_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_110_i2_3_lut_4_lut (.A(n15012), .B(n15001), .C(\array[149] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3249[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_110_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_110_i3_3_lut_4_lut (.A(n15012), .B(n15001), .C(\array[149] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3249[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_110_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_110_i4_3_lut_4_lut (.A(n15012), .B(n15001), .C(\array[149] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3249[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_110_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_110_i5_3_lut_4_lut (.A(n15012), .B(n15001), .C(\array[149] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3249[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_110_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_110_i6_3_lut_4_lut (.A(n15012), .B(n15001), .C(\array[149] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3249[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_110_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_110_i7_3_lut_4_lut (.A(n15012), .B(n15001), .C(\array[149] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3249[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_110_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_110_i8_3_lut_4_lut (.A(n15012), .B(n15001), .C(\array[149] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3249[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_110_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_109_i1_3_lut_4_lut (.A(n15013), .B(n15001), .C(\array[150] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3257[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_109_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_109_i2_3_lut_4_lut (.A(n15013), .B(n15001), .C(\array[150] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3257[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_109_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_109_i3_3_lut_4_lut (.A(n15013), .B(n15001), .C(\array[150] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3257[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_109_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_109_i4_3_lut_4_lut (.A(n15013), .B(n15001), .C(\array[150] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3257[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_109_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_109_i5_3_lut_4_lut (.A(n15013), .B(n15001), .C(\array[150] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3257[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_109_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_109_i6_3_lut_4_lut (.A(n15013), .B(n15001), .C(\array[150] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3257[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_109_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_109_i7_3_lut_4_lut (.A(n15013), .B(n15001), .C(\array[150] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3257[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_109_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_109_i8_3_lut_4_lut (.A(n15013), .B(n15001), .C(\array[150] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3257[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_109_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_108_i1_3_lut_4_lut (.A(n15014), .B(n15001), .C(\array[151] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3265[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_108_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_108_i2_3_lut_4_lut (.A(n15014), .B(n15001), .C(\array[151] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3265[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_108_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_108_i3_3_lut_4_lut (.A(n15014), .B(n15001), .C(\array[151] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3265[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_108_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_108_i4_3_lut_4_lut (.A(n15014), .B(n15001), .C(\array[151] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3265[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_108_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_108_i5_3_lut_4_lut (.A(n15014), .B(n15001), .C(\array[151] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3265[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_108_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_108_i6_3_lut_4_lut (.A(n15014), .B(n15001), .C(\array[151] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3265[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_108_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_108_i7_3_lut_4_lut (.A(n15014), .B(n15001), .C(\array[151] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3265[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_108_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_108_i8_3_lut_4_lut (.A(n15014), .B(n15001), .C(\array[151] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3265[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_108_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_107_i1_3_lut_4_lut (.A(n15015), .B(n15001), .C(\array[152] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3273[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_107_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_107_i2_3_lut_4_lut (.A(n15015), .B(n15001), .C(\array[152] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3273[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_107_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_107_i3_3_lut_4_lut (.A(n15015), .B(n15001), .C(\array[152] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3273[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_107_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_107_i4_3_lut_4_lut (.A(n15015), .B(n15001), .C(\array[152] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3273[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_107_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_107_i5_3_lut_4_lut (.A(n15015), .B(n15001), .C(\array[152] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3273[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_107_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_107_i6_3_lut_4_lut (.A(n15015), .B(n15001), .C(\array[152] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3273[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_107_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_107_i7_3_lut_4_lut (.A(n15015), .B(n15001), .C(\array[152] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3273[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_107_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_107_i8_3_lut_4_lut (.A(n15015), .B(n15001), .C(\array[152] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3273[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_107_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_106_i1_3_lut_4_lut (.A(n15016), .B(n15001), .C(\array[153] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3281[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_106_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_106_i2_3_lut_4_lut (.A(n15016), .B(n15001), .C(\array[153] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3281[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_106_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_106_i3_3_lut_4_lut (.A(n15016), .B(n15001), .C(\array[153] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3281[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_106_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_106_i4_3_lut_4_lut (.A(n15016), .B(n15001), .C(\array[153] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3281[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_106_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_106_i5_3_lut_4_lut (.A(n15016), .B(n15001), .C(\array[153] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3281[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_106_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_106_i6_3_lut_4_lut (.A(n15016), .B(n15001), .C(\array[153] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3281[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_106_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_106_i7_3_lut_4_lut (.A(n15016), .B(n15001), .C(\array[153] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3281[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_106_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_106_i8_3_lut_4_lut (.A(n15016), .B(n15001), .C(\array[153] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3281[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_106_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_105_i1_3_lut_4_lut (.A(n15017), .B(n15001), .C(\array[154] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3289[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_105_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_105_i2_3_lut_4_lut (.A(n15017), .B(n15001), .C(\array[154] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3289[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_105_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_105_i3_3_lut_4_lut (.A(n15017), .B(n15001), .C(\array[154] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3289[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_105_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_105_i4_3_lut_4_lut (.A(n15017), .B(n15001), .C(\array[154] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3289[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_105_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_105_i5_3_lut_4_lut (.A(n15017), .B(n15001), .C(\array[154] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3289[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_105_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_105_i6_3_lut_4_lut (.A(n15017), .B(n15001), .C(\array[154] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3289[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_105_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_105_i7_3_lut_4_lut (.A(n15017), .B(n15001), .C(\array[154] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3289[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_105_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_105_i8_3_lut_4_lut (.A(n15017), .B(n15001), .C(\array[154] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3289[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_105_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_104_i1_3_lut_4_lut (.A(n15018), .B(n15001), .C(\array[155] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3297[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_104_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_104_i2_3_lut_4_lut (.A(n15018), .B(n15001), .C(\array[155] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3297[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_104_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_104_i3_3_lut_4_lut (.A(n15018), .B(n15001), .C(\array[155] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3297[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_104_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_104_i4_3_lut_4_lut (.A(n15018), .B(n15001), .C(\array[155] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3297[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_104_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_104_i5_3_lut_4_lut (.A(n15018), .B(n15001), .C(\array[155] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3297[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_104_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_104_i6_3_lut_4_lut (.A(n15018), .B(n15001), .C(\array[155] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3297[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_104_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_104_i7_3_lut_4_lut (.A(n15018), .B(n15001), .C(\array[155] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3297[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_104_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_104_i8_3_lut_4_lut (.A(n15018), .B(n15001), .C(\array[155] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3297[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_104_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_103_i1_3_lut_4_lut (.A(n15019), .B(n15001), .C(\array[156] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3305[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_103_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_103_i2_3_lut_4_lut (.A(n15019), .B(n15001), .C(\array[156] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3305[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_103_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_103_i3_3_lut_4_lut (.A(n15019), .B(n15001), .C(\array[156] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3305[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_103_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_103_i4_3_lut_4_lut (.A(n15019), .B(n15001), .C(\array[156] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3305[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_103_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_103_i5_3_lut_4_lut (.A(n15019), .B(n15001), .C(\array[156] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3305[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_103_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_103_i6_3_lut_4_lut (.A(n15019), .B(n15001), .C(\array[156] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3305[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_103_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_103_i7_3_lut_4_lut (.A(n15019), .B(n15001), .C(\array[156] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3305[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_103_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_103_i8_3_lut_4_lut (.A(n15019), .B(n15001), .C(\array[156] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3305[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_103_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_102_i1_3_lut_4_lut (.A(n15020), .B(n15001), .C(\array[157] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3313[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_102_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_102_i2_3_lut_4_lut (.A(n15020), .B(n15001), .C(\array[157] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3313[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_102_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_102_i3_3_lut_4_lut (.A(n15020), .B(n15001), .C(\array[157] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3313[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_102_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_102_i4_3_lut_4_lut (.A(n15020), .B(n15001), .C(\array[157] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3313[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_102_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_102_i5_3_lut_4_lut (.A(n15020), .B(n15001), .C(\array[157] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3313[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_102_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_102_i6_3_lut_4_lut (.A(n15020), .B(n15001), .C(\array[157] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3313[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_102_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_102_i7_3_lut_4_lut (.A(n15020), .B(n15001), .C(\array[157] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3313[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_102_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_102_i8_3_lut_4_lut (.A(n15020), .B(n15001), .C(\array[157] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3313[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_102_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_101_i1_3_lut_4_lut (.A(n15021), .B(n15001), .C(\array[158] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3321[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_101_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_101_i2_3_lut_4_lut (.A(n15021), .B(n15001), .C(\array[158] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3321[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_101_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_101_i3_3_lut_4_lut (.A(n15021), .B(n15001), .C(\array[158] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3321[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_101_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_101_i4_3_lut_4_lut (.A(n15021), .B(n15001), .C(\array[158] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3321[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_101_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_101_i5_3_lut_4_lut (.A(n15021), .B(n15001), .C(\array[158] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3321[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_101_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_101_i6_3_lut_4_lut (.A(n15021), .B(n15001), .C(\array[158] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3321[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_101_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_101_i7_3_lut_4_lut (.A(n15021), .B(n15001), .C(\array[158] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3321[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_101_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_101_i8_3_lut_4_lut (.A(n15021), .B(n15001), .C(\array[158] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3321[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_101_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_100_i1_3_lut_4_lut (.A(n15023), .B(n15001), .C(\array[159] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3329[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_100_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_100_i2_3_lut_4_lut (.A(n15023), .B(n15001), .C(\array[159] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3329[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_100_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_100_i3_3_lut_4_lut (.A(n15023), .B(n15001), .C(\array[159] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3329[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_100_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_100_i4_3_lut_4_lut (.A(n15023), .B(n15001), .C(\array[159] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3329[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_100_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_100_i5_3_lut_4_lut (.A(n15023), .B(n15001), .C(\array[159] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3329[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_100_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_100_i6_3_lut_4_lut (.A(n15023), .B(n15001), .C(\array[159] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3329[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_100_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_100_i7_3_lut_4_lut (.A(n15023), .B(n15001), .C(\array[159] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3329[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_100_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_100_i8_3_lut_4_lut (.A(n15023), .B(n15001), .C(\array[159] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3329[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_100_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_99_i1_3_lut_4_lut (.A(n15007), .B(n15002), .C(\array[160] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3337[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_99_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_99_i2_3_lut_4_lut (.A(n15007), .B(n15002), .C(\array[160] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3337[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_99_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_99_i3_3_lut_4_lut (.A(n15007), .B(n15002), .C(\array[160] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3337[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_99_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_99_i4_3_lut_4_lut (.A(n15007), .B(n15002), .C(\array[160] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3337[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_99_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_99_i5_3_lut_4_lut (.A(n15007), .B(n15002), .C(\array[160] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3337[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_99_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_99_i6_3_lut_4_lut (.A(n15007), .B(n15002), .C(\array[160] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3337[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_99_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_99_i7_3_lut_4_lut (.A(n15007), .B(n15002), .C(\array[160] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3337[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_99_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_99_i8_3_lut_4_lut (.A(n15007), .B(n15002), .C(\array[160] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3337[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_99_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_98_i1_3_lut_4_lut (.A(n15008), .B(n15002), .C(\array[161] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3345[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_98_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_98_i2_3_lut_4_lut (.A(n15008), .B(n15002), .C(\array[161] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3345[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_98_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_98_i3_3_lut_4_lut (.A(n15008), .B(n15002), .C(\array[161] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3345[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_98_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_98_i4_3_lut_4_lut (.A(n15008), .B(n15002), .C(\array[161] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3345[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_98_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_98_i5_3_lut_4_lut (.A(n15008), .B(n15002), .C(\array[161] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3345[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_98_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_98_i6_3_lut_4_lut (.A(n15008), .B(n15002), .C(\array[161] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3345[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_98_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_98_i7_3_lut_4_lut (.A(n15008), .B(n15002), .C(\array[161] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3345[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_98_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_98_i8_3_lut_4_lut (.A(n15008), .B(n15002), .C(\array[161] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3345[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_98_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_97_i1_3_lut_4_lut (.A(n15009), .B(n15002), .C(\array[162] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3353[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_97_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_97_i2_3_lut_4_lut (.A(n15009), .B(n15002), .C(\array[162] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3353[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_97_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_97_i3_3_lut_4_lut (.A(n15009), .B(n15002), .C(\array[162] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3353[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_97_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_97_i4_3_lut_4_lut (.A(n15009), .B(n15002), .C(\array[162] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3353[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_97_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_97_i5_3_lut_4_lut (.A(n15009), .B(n15002), .C(\array[162] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3353[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_97_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_97_i6_3_lut_4_lut (.A(n15009), .B(n15002), .C(\array[162] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3353[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_97_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_97_i7_3_lut_4_lut (.A(n15009), .B(n15002), .C(\array[162] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3353[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_97_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_97_i8_3_lut_4_lut (.A(n15009), .B(n15002), .C(\array[162] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3353[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_97_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_96_i1_3_lut_4_lut (.A(n15010), .B(n15002), .C(\array[163] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3361[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_96_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_96_i2_3_lut_4_lut (.A(n15010), .B(n15002), .C(\array[163] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3361[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_96_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_96_i3_3_lut_4_lut (.A(n15010), .B(n15002), .C(\array[163] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3361[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_96_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_96_i4_3_lut_4_lut (.A(n15010), .B(n15002), .C(\array[163] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3361[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_96_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_96_i5_3_lut_4_lut (.A(n15010), .B(n15002), .C(\array[163] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3361[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_96_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_96_i6_3_lut_4_lut (.A(n15010), .B(n15002), .C(\array[163] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3361[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_96_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_96_i7_3_lut_4_lut (.A(n15010), .B(n15002), .C(\array[163] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3361[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_96_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_96_i8_3_lut_4_lut (.A(n15010), .B(n15002), .C(\array[163] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3361[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_96_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_95_i1_3_lut_4_lut (.A(n15011), .B(n15002), .C(\array[164] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3369[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_95_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_95_i2_3_lut_4_lut (.A(n15011), .B(n15002), .C(\array[164] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3369[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_95_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_95_i3_3_lut_4_lut (.A(n15011), .B(n15002), .C(\array[164] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3369[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_95_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_95_i4_3_lut_4_lut (.A(n15011), .B(n15002), .C(\array[164] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3369[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_95_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_95_i5_3_lut_4_lut (.A(n15011), .B(n15002), .C(\array[164] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3369[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_95_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_95_i6_3_lut_4_lut (.A(n15011), .B(n15002), .C(\array[164] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3369[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_95_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_95_i7_3_lut_4_lut (.A(n15011), .B(n15002), .C(\array[164] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3369[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_95_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_95_i8_3_lut_4_lut (.A(n15011), .B(n15002), .C(\array[164] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3369[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_95_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_94_i1_3_lut_4_lut (.A(n15012), .B(n15002), .C(\array[165] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3377[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_94_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_94_i2_3_lut_4_lut (.A(n15012), .B(n15002), .C(\array[165] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3377[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_94_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_94_i3_3_lut_4_lut (.A(n15012), .B(n15002), .C(\array[165] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3377[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_94_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_94_i4_3_lut_4_lut (.A(n15012), .B(n15002), .C(\array[165] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3377[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_94_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_94_i5_3_lut_4_lut (.A(n15012), .B(n15002), .C(\array[165] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3377[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_94_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_94_i6_3_lut_4_lut (.A(n15012), .B(n15002), .C(\array[165] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3377[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_94_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_94_i7_3_lut_4_lut (.A(n15012), .B(n15002), .C(\array[165] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3377[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_94_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_94_i8_3_lut_4_lut (.A(n15012), .B(n15002), .C(\array[165] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3377[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_94_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_93_i1_3_lut_4_lut (.A(n15013), .B(n15002), .C(\array[166] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3385[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_93_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_93_i2_3_lut_4_lut (.A(n15013), .B(n15002), .C(\array[166] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3385[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_93_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_93_i3_3_lut_4_lut (.A(n15013), .B(n15002), .C(\array[166] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3385[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_93_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_93_i4_3_lut_4_lut (.A(n15013), .B(n15002), .C(\array[166] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3385[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_93_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_93_i5_3_lut_4_lut (.A(n15013), .B(n15002), .C(\array[166] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3385[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_93_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_93_i6_3_lut_4_lut (.A(n15013), .B(n15002), .C(\array[166] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3385[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_93_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_93_i7_3_lut_4_lut (.A(n15013), .B(n15002), .C(\array[166] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3385[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_93_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_93_i8_3_lut_4_lut (.A(n15013), .B(n15002), .C(\array[166] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3385[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_93_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_92_i1_3_lut_4_lut (.A(n15014), .B(n15002), .C(\array[167] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3393[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_92_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_92_i2_3_lut_4_lut (.A(n15014), .B(n15002), .C(\array[167] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3393[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_92_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_92_i3_3_lut_4_lut (.A(n15014), .B(n15002), .C(\array[167] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3393[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_92_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_92_i4_3_lut_4_lut (.A(n15014), .B(n15002), .C(\array[167] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3393[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_92_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_92_i5_3_lut_4_lut (.A(n15014), .B(n15002), .C(\array[167] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3393[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_92_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_92_i6_3_lut_4_lut (.A(n15014), .B(n15002), .C(\array[167] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3393[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_92_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_92_i7_3_lut_4_lut (.A(n15014), .B(n15002), .C(\array[167] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3393[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_92_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_92_i8_3_lut_4_lut (.A(n15014), .B(n15002), .C(\array[167] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3393[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_92_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_91_i1_3_lut_4_lut (.A(n15015), .B(n15002), .C(\array[168] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3401[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_91_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_91_i2_3_lut_4_lut (.A(n15015), .B(n15002), .C(\array[168] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3401[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_91_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_91_i3_3_lut_4_lut (.A(n15015), .B(n15002), .C(\array[168] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3401[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_91_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_91_i4_3_lut_4_lut (.A(n15015), .B(n15002), .C(\array[168] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3401[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_91_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_91_i5_3_lut_4_lut (.A(n15015), .B(n15002), .C(\array[168] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3401[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_91_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_91_i6_3_lut_4_lut (.A(n15015), .B(n15002), .C(\array[168] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3401[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_91_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_91_i7_3_lut_4_lut (.A(n15015), .B(n15002), .C(\array[168] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3401[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_91_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_91_i8_3_lut_4_lut (.A(n15015), .B(n15002), .C(\array[168] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3401[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_91_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_90_i1_3_lut_4_lut (.A(n15016), .B(n15002), .C(\array[169] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3409[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_90_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_90_i2_3_lut_4_lut (.A(n15016), .B(n15002), .C(\array[169] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3409[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_90_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_90_i3_3_lut_4_lut (.A(n15016), .B(n15002), .C(\array[169] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3409[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_90_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_90_i4_3_lut_4_lut (.A(n15016), .B(n15002), .C(\array[169] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3409[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_90_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_90_i5_3_lut_4_lut (.A(n15016), .B(n15002), .C(\array[169] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3409[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_90_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_90_i6_3_lut_4_lut (.A(n15016), .B(n15002), .C(\array[169] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3409[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_90_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_90_i7_3_lut_4_lut (.A(n15016), .B(n15002), .C(\array[169] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3409[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_90_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_90_i8_3_lut_4_lut (.A(n15016), .B(n15002), .C(\array[169] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3409[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_90_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_89_i1_3_lut_4_lut (.A(n15017), .B(n15002), .C(\array[170] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3417[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_89_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_89_i2_3_lut_4_lut (.A(n15017), .B(n15002), .C(\array[170] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3417[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_89_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_89_i3_3_lut_4_lut (.A(n15017), .B(n15002), .C(\array[170] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3417[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_89_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_89_i4_3_lut_4_lut (.A(n15017), .B(n15002), .C(\array[170] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3417[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_89_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_89_i5_3_lut_4_lut (.A(n15017), .B(n15002), .C(\array[170] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3417[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_89_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_89_i6_3_lut_4_lut (.A(n15017), .B(n15002), .C(\array[170] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3417[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_89_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_89_i7_3_lut_4_lut (.A(n15017), .B(n15002), .C(\array[170] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3417[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_89_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_89_i8_3_lut_4_lut (.A(n15017), .B(n15002), .C(\array[170] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3417[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_89_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_88_i1_3_lut_4_lut (.A(n15018), .B(n15002), .C(\array[171] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3425[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_88_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_88_i2_3_lut_4_lut (.A(n15018), .B(n15002), .C(\array[171] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3425[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_88_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_88_i3_3_lut_4_lut (.A(n15018), .B(n15002), .C(\array[171] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3425[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_88_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_88_i4_3_lut_4_lut (.A(n15018), .B(n15002), .C(\array[171] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3425[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_88_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_88_i5_3_lut_4_lut (.A(n15018), .B(n15002), .C(\array[171] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3425[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_88_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_88_i6_3_lut_4_lut (.A(n15018), .B(n15002), .C(\array[171] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3425[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_88_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_88_i7_3_lut_4_lut (.A(n15018), .B(n15002), .C(\array[171] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3425[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_88_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_88_i8_3_lut_4_lut (.A(n15018), .B(n15002), .C(\array[171] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3425[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_88_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_87_i1_3_lut_4_lut (.A(n15019), .B(n15002), .C(\array[172] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3433[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_87_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_87_i2_3_lut_4_lut (.A(n15019), .B(n15002), .C(\array[172] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3433[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_87_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_87_i3_3_lut_4_lut (.A(n15019), .B(n15002), .C(\array[172] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3433[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_87_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_87_i4_3_lut_4_lut (.A(n15019), .B(n15002), .C(\array[172] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3433[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_87_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_87_i5_3_lut_4_lut (.A(n15019), .B(n15002), .C(\array[172] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3433[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_87_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_87_i6_3_lut_4_lut (.A(n15019), .B(n15002), .C(\array[172] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3433[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_87_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_87_i7_3_lut_4_lut (.A(n15019), .B(n15002), .C(\array[172] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3433[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_87_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_87_i8_3_lut_4_lut (.A(n15019), .B(n15002), .C(\array[172] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3433[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_87_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_86_i1_3_lut_4_lut (.A(n15020), .B(n15002), .C(\array[173] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3441[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_86_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_86_i2_3_lut_4_lut (.A(n15020), .B(n15002), .C(\array[173] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3441[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_86_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_86_i3_3_lut_4_lut (.A(n15020), .B(n15002), .C(\array[173] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3441[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_86_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_86_i4_3_lut_4_lut (.A(n15020), .B(n15002), .C(\array[173] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3441[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_86_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_86_i5_3_lut_4_lut (.A(n15020), .B(n15002), .C(\array[173] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3441[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_86_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_86_i6_3_lut_4_lut (.A(n15020), .B(n15002), .C(\array[173] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3441[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_86_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_86_i7_3_lut_4_lut (.A(n15020), .B(n15002), .C(\array[173] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3441[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_86_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_86_i8_3_lut_4_lut (.A(n15020), .B(n15002), .C(\array[173] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3441[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_86_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i1_3_lut_4_lut (.A(n15021), .B(n15002), .C(\array[174] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3449[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_85_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i2_3_lut_4_lut (.A(n15021), .B(n15002), .C(\array[174] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3449[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_85_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i3_3_lut_4_lut (.A(n15021), .B(n15002), .C(\array[174] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3449[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_85_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i4_3_lut_4_lut (.A(n15021), .B(n15002), .C(\array[174] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3449[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_85_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i5_3_lut_4_lut (.A(n15021), .B(n15002), .C(\array[174] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3449[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_85_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i6_3_lut_4_lut (.A(n15021), .B(n15002), .C(\array[174] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3449[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_85_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i7_3_lut_4_lut (.A(n15021), .B(n15002), .C(\array[174] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3449[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_85_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_85_i8_3_lut_4_lut (.A(n15021), .B(n15002), .C(\array[174] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3449[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_85_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_84_i1_3_lut_4_lut (.A(n15023), .B(n15002), .C(\array[175] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3457[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_84_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_84_i2_3_lut_4_lut (.A(n15023), .B(n15002), .C(\array[175] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3457[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_84_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_84_i3_3_lut_4_lut (.A(n15023), .B(n15002), .C(\array[175] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3457[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_84_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_84_i4_3_lut_4_lut (.A(n15023), .B(n15002), .C(\array[175] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3457[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_84_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_84_i5_3_lut_4_lut (.A(n15023), .B(n15002), .C(\array[175] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3457[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_84_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_84_i6_3_lut_4_lut (.A(n15023), .B(n15002), .C(\array[175] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3457[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_84_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_84_i7_3_lut_4_lut (.A(n15023), .B(n15002), .C(\array[175] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3457[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_84_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_84_i8_3_lut_4_lut (.A(n15023), .B(n15002), .C(\array[175] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3457[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_84_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_83_i1_3_lut_4_lut (.A(n15007), .B(n15003), .C(\array[176] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3465[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_83_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_83_i2_3_lut_4_lut (.A(n15007), .B(n15003), .C(\array[176] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3465[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_83_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_83_i3_3_lut_4_lut (.A(n15007), .B(n15003), .C(\array[176] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3465[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_83_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_83_i4_3_lut_4_lut (.A(n15007), .B(n15003), .C(\array[176] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3465[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_83_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_83_i5_3_lut_4_lut (.A(n15007), .B(n15003), .C(\array[176] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3465[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_83_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_83_i6_3_lut_4_lut (.A(n15007), .B(n15003), .C(\array[176] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3465[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_83_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_83_i7_3_lut_4_lut (.A(n15007), .B(n15003), .C(\array[176] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3465[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_83_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_83_i8_3_lut_4_lut (.A(n15007), .B(n15003), .C(\array[176] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3465[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_83_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_82_i1_3_lut_4_lut (.A(n15008), .B(n15003), .C(\array[177] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3473[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_82_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_82_i2_3_lut_4_lut (.A(n15008), .B(n15003), .C(\array[177] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3473[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_82_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_82_i3_3_lut_4_lut (.A(n15008), .B(n15003), .C(\array[177] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3473[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_82_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_82_i4_3_lut_4_lut (.A(n15008), .B(n15003), .C(\array[177] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3473[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_82_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_82_i5_3_lut_4_lut (.A(n15008), .B(n15003), .C(\array[177] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3473[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_82_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_82_i6_3_lut_4_lut (.A(n15008), .B(n15003), .C(\array[177] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3473[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_82_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_82_i7_3_lut_4_lut (.A(n15008), .B(n15003), .C(\array[177] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3473[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_82_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_82_i8_3_lut_4_lut (.A(n15008), .B(n15003), .C(\array[177] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3473[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_82_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_81_i1_3_lut_4_lut (.A(n15009), .B(n15003), .C(\array[178] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3481[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_81_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_81_i2_3_lut_4_lut (.A(n15009), .B(n15003), .C(\array[178] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3481[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_81_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_81_i3_3_lut_4_lut (.A(n15009), .B(n15003), .C(\array[178] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3481[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_81_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_81_i4_3_lut_4_lut (.A(n15009), .B(n15003), .C(\array[178] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3481[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_81_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_81_i5_3_lut_4_lut (.A(n15009), .B(n15003), .C(\array[178] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3481[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_81_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_81_i6_3_lut_4_lut (.A(n15009), .B(n15003), .C(\array[178] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3481[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_81_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_81_i7_3_lut_4_lut (.A(n15009), .B(n15003), .C(\array[178] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3481[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_81_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_81_i8_3_lut_4_lut (.A(n15009), .B(n15003), .C(\array[178] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3481[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_81_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_80_i1_3_lut_4_lut (.A(n15010), .B(n15003), .C(\array[179] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3489[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_80_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_80_i2_3_lut_4_lut (.A(n15010), .B(n15003), .C(\array[179] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3489[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_80_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_80_i3_3_lut_4_lut (.A(n15010), .B(n15003), .C(\array[179] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3489[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_80_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_80_i4_3_lut_4_lut (.A(n15010), .B(n15003), .C(\array[179] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3489[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_80_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_80_i5_3_lut_4_lut (.A(n15010), .B(n15003), .C(\array[179] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3489[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_80_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_80_i6_3_lut_4_lut (.A(n15010), .B(n15003), .C(\array[179] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3489[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_80_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_80_i7_3_lut_4_lut (.A(n15010), .B(n15003), .C(\array[179] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3489[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_80_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_80_i8_3_lut_4_lut (.A(n15010), .B(n15003), .C(\array[179] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3489[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_80_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_79_i1_3_lut_4_lut (.A(n15011), .B(n15003), .C(\array[180] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3497[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_79_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_79_i2_3_lut_4_lut (.A(n15011), .B(n15003), .C(\array[180] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3497[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_79_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_79_i3_3_lut_4_lut (.A(n15011), .B(n15003), .C(\array[180] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3497[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_79_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_79_i4_3_lut_4_lut (.A(n15011), .B(n15003), .C(\array[180] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3497[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_79_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_79_i5_3_lut_4_lut (.A(n15011), .B(n15003), .C(\array[180] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3497[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_79_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_79_i6_3_lut_4_lut (.A(n15011), .B(n15003), .C(\array[180] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3497[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_79_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_79_i7_3_lut_4_lut (.A(n15011), .B(n15003), .C(\array[180] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3497[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_79_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_79_i8_3_lut_4_lut (.A(n15011), .B(n15003), .C(\array[180] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3497[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_79_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_78_i1_3_lut_4_lut (.A(n15012), .B(n15003), .C(\array[181] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3505[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_78_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_78_i2_3_lut_4_lut (.A(n15012), .B(n15003), .C(\array[181] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3505[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_78_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_78_i3_3_lut_4_lut (.A(n15012), .B(n15003), .C(\array[181] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3505[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_78_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_78_i4_3_lut_4_lut (.A(n15012), .B(n15003), .C(\array[181] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3505[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_78_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_78_i5_3_lut_4_lut (.A(n15012), .B(n15003), .C(\array[181] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3505[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_78_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_78_i6_3_lut_4_lut (.A(n15012), .B(n15003), .C(\array[181] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3505[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_78_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_78_i7_3_lut_4_lut (.A(n15012), .B(n15003), .C(\array[181] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3505[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_78_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_78_i8_3_lut_4_lut (.A(n15012), .B(n15003), .C(\array[181] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3505[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_78_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_77_i1_3_lut_4_lut (.A(n15013), .B(n15003), .C(\array[182] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3513[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_77_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_77_i2_3_lut_4_lut (.A(n15013), .B(n15003), .C(\array[182] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3513[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_77_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_77_i3_3_lut_4_lut (.A(n15013), .B(n15003), .C(\array[182] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3513[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_77_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_77_i4_3_lut_4_lut (.A(n15013), .B(n15003), .C(\array[182] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3513[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_77_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_77_i5_3_lut_4_lut (.A(n15013), .B(n15003), .C(\array[182] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3513[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_77_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_77_i6_3_lut_4_lut (.A(n15013), .B(n15003), .C(\array[182] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3513[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_77_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_77_i7_3_lut_4_lut (.A(n15013), .B(n15003), .C(\array[182] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3513[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_77_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_77_i8_3_lut_4_lut (.A(n15013), .B(n15003), .C(\array[182] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3513[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_77_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_76_i1_3_lut_4_lut (.A(n15014), .B(n15003), .C(\array[183] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3521[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_76_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_76_i2_3_lut_4_lut (.A(n15014), .B(n15003), .C(\array[183] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3521[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_76_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_76_i3_3_lut_4_lut (.A(n15014), .B(n15003), .C(\array[183] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3521[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_76_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_76_i4_3_lut_4_lut (.A(n15014), .B(n15003), .C(\array[183] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3521[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_76_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_76_i5_3_lut_4_lut (.A(n15014), .B(n15003), .C(\array[183] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3521[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_76_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_76_i6_3_lut_4_lut (.A(n15014), .B(n15003), .C(\array[183] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3521[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_76_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_76_i7_3_lut_4_lut (.A(n15014), .B(n15003), .C(\array[183] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3521[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_76_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_76_i8_3_lut_4_lut (.A(n15014), .B(n15003), .C(\array[183] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3521[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_76_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_75_i1_3_lut_4_lut (.A(n15015), .B(n15003), .C(\array[184] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3529[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_75_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_75_i2_3_lut_4_lut (.A(n15015), .B(n15003), .C(\array[184] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3529[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_75_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_75_i3_3_lut_4_lut (.A(n15015), .B(n15003), .C(\array[184] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3529[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_75_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_75_i4_3_lut_4_lut (.A(n15015), .B(n15003), .C(\array[184] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3529[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_75_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_75_i5_3_lut_4_lut (.A(n15015), .B(n15003), .C(\array[184] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3529[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_75_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_75_i6_3_lut_4_lut (.A(n15015), .B(n15003), .C(\array[184] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3529[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_75_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_75_i7_3_lut_4_lut (.A(n15015), .B(n15003), .C(\array[184] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3529[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_75_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_75_i8_3_lut_4_lut (.A(n15015), .B(n15003), .C(\array[184] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3529[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_75_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_74_i1_3_lut_4_lut (.A(n15016), .B(n15003), .C(\array[185] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3537[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_74_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_74_i2_3_lut_4_lut (.A(n15016), .B(n15003), .C(\array[185] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3537[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_74_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_74_i3_3_lut_4_lut (.A(n15016), .B(n15003), .C(\array[185] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3537[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_74_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_74_i4_3_lut_4_lut (.A(n15016), .B(n15003), .C(\array[185] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3537[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_74_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_74_i5_3_lut_4_lut (.A(n15016), .B(n15003), .C(\array[185] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3537[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_74_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_74_i6_3_lut_4_lut (.A(n15016), .B(n15003), .C(\array[185] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3537[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_74_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_74_i7_3_lut_4_lut (.A(n15016), .B(n15003), .C(\array[185] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3537[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_74_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_74_i8_3_lut_4_lut (.A(n15016), .B(n15003), .C(\array[185] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3537[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_74_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_73_i1_3_lut_4_lut (.A(n15017), .B(n15003), .C(\array[186] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3545[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_73_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_73_i2_3_lut_4_lut (.A(n15017), .B(n15003), .C(\array[186] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3545[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_73_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_73_i3_3_lut_4_lut (.A(n15017), .B(n15003), .C(\array[186] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3545[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_73_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_73_i4_3_lut_4_lut (.A(n15017), .B(n15003), .C(\array[186] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3545[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_73_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_73_i5_3_lut_4_lut (.A(n15017), .B(n15003), .C(\array[186] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3545[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_73_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_73_i6_3_lut_4_lut (.A(n15017), .B(n15003), .C(\array[186] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3545[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_73_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_73_i7_3_lut_4_lut (.A(n15017), .B(n15003), .C(\array[186] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3545[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_73_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_73_i8_3_lut_4_lut (.A(n15017), .B(n15003), .C(\array[186] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3545[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_73_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_72_i1_3_lut_4_lut (.A(n15018), .B(n15003), .C(\array[187] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3553[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_72_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_72_i2_3_lut_4_lut (.A(n15018), .B(n15003), .C(\array[187] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3553[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_72_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_72_i3_3_lut_4_lut (.A(n15018), .B(n15003), .C(\array[187] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3553[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_72_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_72_i4_3_lut_4_lut (.A(n15018), .B(n15003), .C(\array[187] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3553[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_72_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_72_i5_3_lut_4_lut (.A(n15018), .B(n15003), .C(\array[187] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3553[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_72_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_72_i6_3_lut_4_lut (.A(n15018), .B(n15003), .C(\array[187] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3553[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_72_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_72_i7_3_lut_4_lut (.A(n15018), .B(n15003), .C(\array[187] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3553[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_72_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_72_i8_3_lut_4_lut (.A(n15018), .B(n15003), .C(\array[187] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3553[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_72_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_71_i1_3_lut_4_lut (.A(n15019), .B(n15003), .C(\array[188] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3561[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_71_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_71_i2_3_lut_4_lut (.A(n15019), .B(n15003), .C(\array[188] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3561[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_71_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_71_i3_3_lut_4_lut (.A(n15019), .B(n15003), .C(\array[188] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3561[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_71_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_71_i4_3_lut_4_lut (.A(n15019), .B(n15003), .C(\array[188] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3561[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_71_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_71_i5_3_lut_4_lut (.A(n15019), .B(n15003), .C(\array[188] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3561[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_71_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_71_i6_3_lut_4_lut (.A(n15019), .B(n15003), .C(\array[188] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3561[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_71_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_71_i7_3_lut_4_lut (.A(n15019), .B(n15003), .C(\array[188] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3561[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_71_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_71_i8_3_lut_4_lut (.A(n15019), .B(n15003), .C(\array[188] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3561[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_71_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_70_i1_3_lut_4_lut (.A(n15020), .B(n15003), .C(\array[189] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3569[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_70_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_70_i2_3_lut_4_lut (.A(n15020), .B(n15003), .C(\array[189] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3569[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_70_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_70_i3_3_lut_4_lut (.A(n15020), .B(n15003), .C(\array[189] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3569[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_70_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_70_i4_3_lut_4_lut (.A(n15020), .B(n15003), .C(\array[189] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3569[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_70_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_70_i5_3_lut_4_lut (.A(n15020), .B(n15003), .C(\array[189] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3569[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_70_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_70_i6_3_lut_4_lut (.A(n15020), .B(n15003), .C(\array[189] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3569[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_70_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_70_i7_3_lut_4_lut (.A(n15020), .B(n15003), .C(\array[189] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3569[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_70_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_70_i8_3_lut_4_lut (.A(n15020), .B(n15003), .C(\array[189] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3569[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_70_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_69_i1_3_lut_4_lut (.A(n15021), .B(n15003), .C(\array[190] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3577[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_69_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_69_i2_3_lut_4_lut (.A(n15021), .B(n15003), .C(\array[190] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3577[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_69_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_69_i3_3_lut_4_lut (.A(n15021), .B(n15003), .C(\array[190] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3577[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_69_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_69_i4_3_lut_4_lut (.A(n15021), .B(n15003), .C(\array[190] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3577[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_69_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_69_i5_3_lut_4_lut (.A(n15021), .B(n15003), .C(\array[190] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3577[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_69_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_69_i6_3_lut_4_lut (.A(n15021), .B(n15003), .C(\array[190] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3577[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_69_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_69_i7_3_lut_4_lut (.A(n15021), .B(n15003), .C(\array[190] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3577[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_69_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_69_i8_3_lut_4_lut (.A(n15021), .B(n15003), .C(\array[190] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3577[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_69_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_68_i1_3_lut_4_lut (.A(n15023), .B(n15003), .C(\array[191] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3585[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_68_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_68_i2_3_lut_4_lut (.A(n15023), .B(n15003), .C(\array[191] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3585[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_68_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_68_i3_3_lut_4_lut (.A(n15023), .B(n15003), .C(\array[191] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3585[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_68_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_68_i4_3_lut_4_lut (.A(n15023), .B(n15003), .C(\array[191] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3585[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_68_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_68_i5_3_lut_4_lut (.A(n15023), .B(n15003), .C(\array[191] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3585[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_68_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_68_i6_3_lut_4_lut (.A(n15023), .B(n15003), .C(\array[191] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3585[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_68_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_68_i7_3_lut_4_lut (.A(n15023), .B(n15003), .C(\array[191] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3585[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_68_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_68_i8_3_lut_4_lut (.A(n15023), .B(n15003), .C(\array[191] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3585[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_68_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_67_i1_3_lut_4_lut (.A(n15007), .B(n15004), .C(\array[192] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3593[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_67_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_67_i2_3_lut_4_lut (.A(n15007), .B(n15004), .C(\array[192] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3593[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_67_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_67_i3_3_lut_4_lut (.A(n15007), .B(n15004), .C(\array[192] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3593[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_67_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_67_i4_3_lut_4_lut (.A(n15007), .B(n15004), .C(\array[192] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3593[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_67_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_67_i5_3_lut_4_lut (.A(n15007), .B(n15004), .C(\array[192] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3593[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_67_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_67_i6_3_lut_4_lut (.A(n15007), .B(n15004), .C(\array[192] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3593[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_67_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_67_i7_3_lut_4_lut (.A(n15007), .B(n15004), .C(\array[192] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3593[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_67_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_67_i8_3_lut_4_lut (.A(n15007), .B(n15004), .C(\array[192] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3593[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_67_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_66_i1_3_lut_4_lut (.A(n15008), .B(n15004), .C(\array[193] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3601[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_66_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_66_i2_3_lut_4_lut (.A(n15008), .B(n15004), .C(\array[193] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3601[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_66_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_66_i3_3_lut_4_lut (.A(n15008), .B(n15004), .C(\array[193] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3601[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_66_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_66_i4_3_lut_4_lut (.A(n15008), .B(n15004), .C(\array[193] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3601[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_66_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_66_i5_3_lut_4_lut (.A(n15008), .B(n15004), .C(\array[193] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3601[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_66_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_66_i6_3_lut_4_lut (.A(n15008), .B(n15004), .C(\array[193] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3601[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_66_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_66_i7_3_lut_4_lut (.A(n15008), .B(n15004), .C(\array[193] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3601[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_66_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_66_i8_3_lut_4_lut (.A(n15008), .B(n15004), .C(\array[193] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3601[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_66_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_65_i1_3_lut_4_lut (.A(n15009), .B(n15004), .C(\array[194] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3609[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_65_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_65_i2_3_lut_4_lut (.A(n15009), .B(n15004), .C(\array[194] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3609[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_65_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_65_i3_3_lut_4_lut (.A(n15009), .B(n15004), .C(\array[194] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3609[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_65_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_65_i4_3_lut_4_lut (.A(n15009), .B(n15004), .C(\array[194] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3609[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_65_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_65_i5_3_lut_4_lut (.A(n15009), .B(n15004), .C(\array[194] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3609[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_65_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_65_i6_3_lut_4_lut (.A(n15009), .B(n15004), .C(\array[194] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3609[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_65_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_65_i7_3_lut_4_lut (.A(n15009), .B(n15004), .C(\array[194] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3609[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_65_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_65_i8_3_lut_4_lut (.A(n15009), .B(n15004), .C(\array[194] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3609[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_65_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_64_i1_3_lut_4_lut (.A(n15010), .B(n15004), .C(\array[195] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3617[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_64_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_64_i2_3_lut_4_lut (.A(n15010), .B(n15004), .C(\array[195] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3617[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_64_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_64_i3_3_lut_4_lut (.A(n15010), .B(n15004), .C(\array[195] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3617[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_64_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_64_i4_3_lut_4_lut (.A(n15010), .B(n15004), .C(\array[195] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3617[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_64_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_64_i5_3_lut_4_lut (.A(n15010), .B(n15004), .C(\array[195] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3617[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_64_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_64_i6_3_lut_4_lut (.A(n15010), .B(n15004), .C(\array[195] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3617[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_64_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_64_i7_3_lut_4_lut (.A(n15010), .B(n15004), .C(\array[195] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3617[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_64_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_64_i8_3_lut_4_lut (.A(n15010), .B(n15004), .C(\array[195] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3617[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_64_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_63_i1_3_lut_4_lut (.A(n15011), .B(n15004), .C(\array[196] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3625[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_63_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_63_i2_3_lut_4_lut (.A(n15011), .B(n15004), .C(\array[196] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3625[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_63_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_63_i3_3_lut_4_lut (.A(n15011), .B(n15004), .C(\array[196] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3625[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_63_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_63_i4_3_lut_4_lut (.A(n15011), .B(n15004), .C(\array[196] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3625[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_63_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_63_i5_3_lut_4_lut (.A(n15011), .B(n15004), .C(\array[196] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3625[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_63_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_63_i6_3_lut_4_lut (.A(n15011), .B(n15004), .C(\array[196] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3625[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_63_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_63_i7_3_lut_4_lut (.A(n15011), .B(n15004), .C(\array[196] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3625[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_63_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_63_i8_3_lut_4_lut (.A(n15011), .B(n15004), .C(\array[196] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3625[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_63_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_62_i1_3_lut_4_lut (.A(n15012), .B(n15004), .C(\array[197] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3633[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_62_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_62_i2_3_lut_4_lut (.A(n15012), .B(n15004), .C(\array[197] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3633[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_62_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_62_i3_3_lut_4_lut (.A(n15012), .B(n15004), .C(\array[197] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3633[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_62_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_62_i4_3_lut_4_lut (.A(n15012), .B(n15004), .C(\array[197] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3633[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_62_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_62_i5_3_lut_4_lut (.A(n15012), .B(n15004), .C(\array[197] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3633[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_62_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_62_i6_3_lut_4_lut (.A(n15012), .B(n15004), .C(\array[197] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3633[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_62_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_62_i7_3_lut_4_lut (.A(n15012), .B(n15004), .C(\array[197] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3633[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_62_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_62_i8_3_lut_4_lut (.A(n15012), .B(n15004), .C(\array[197] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3633[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_62_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_61_i1_3_lut_4_lut (.A(n15013), .B(n15004), .C(\array[198] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3641[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_61_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_61_i2_3_lut_4_lut (.A(n15013), .B(n15004), .C(\array[198] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3641[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_61_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_61_i3_3_lut_4_lut (.A(n15013), .B(n15004), .C(\array[198] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3641[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_61_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_61_i4_3_lut_4_lut (.A(n15013), .B(n15004), .C(\array[198] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3641[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_61_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_61_i5_3_lut_4_lut (.A(n15013), .B(n15004), .C(\array[198] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3641[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_61_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_61_i6_3_lut_4_lut (.A(n15013), .B(n15004), .C(\array[198] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3641[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_61_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_61_i7_3_lut_4_lut (.A(n15013), .B(n15004), .C(\array[198] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3641[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_61_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_61_i8_3_lut_4_lut (.A(n15013), .B(n15004), .C(\array[198] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3641[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_61_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_60_i1_3_lut_4_lut (.A(n15014), .B(n15004), .C(\array[199] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3649[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_60_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_60_i2_3_lut_4_lut (.A(n15014), .B(n15004), .C(\array[199] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3649[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_60_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_60_i3_3_lut_4_lut (.A(n15014), .B(n15004), .C(\array[199] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3649[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_60_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_60_i4_3_lut_4_lut (.A(n15014), .B(n15004), .C(\array[199] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3649[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_60_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_60_i5_3_lut_4_lut (.A(n15014), .B(n15004), .C(\array[199] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3649[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_60_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_60_i6_3_lut_4_lut (.A(n15014), .B(n15004), .C(\array[199] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3649[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_60_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_60_i7_3_lut_4_lut (.A(n15014), .B(n15004), .C(\array[199] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3649[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_60_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_60_i8_3_lut_4_lut (.A(n15014), .B(n15004), .C(\array[199] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3649[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_60_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_59_i1_3_lut_4_lut (.A(n15015), .B(n15004), .C(\array[200] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3657[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_59_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_59_i2_3_lut_4_lut (.A(n15015), .B(n15004), .C(\array[200] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3657[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_59_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_59_i3_3_lut_4_lut (.A(n15015), .B(n15004), .C(\array[200] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3657[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_59_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_59_i4_3_lut_4_lut (.A(n15015), .B(n15004), .C(\array[200] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3657[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_59_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_59_i5_3_lut_4_lut (.A(n15015), .B(n15004), .C(\array[200] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3657[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_59_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_59_i6_3_lut_4_lut (.A(n15015), .B(n15004), .C(\array[200] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3657[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_59_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_59_i7_3_lut_4_lut (.A(n15015), .B(n15004), .C(\array[200] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3657[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_59_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_59_i8_3_lut_4_lut (.A(n15015), .B(n15004), .C(\array[200] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3657[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_59_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_58_i1_3_lut_4_lut (.A(n15016), .B(n15004), .C(\array[201] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3665[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_58_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_58_i2_3_lut_4_lut (.A(n15016), .B(n15004), .C(\array[201] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3665[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_58_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_58_i3_3_lut_4_lut (.A(n15016), .B(n15004), .C(\array[201] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3665[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_58_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_58_i4_3_lut_4_lut (.A(n15016), .B(n15004), .C(\array[201] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3665[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_58_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_58_i5_3_lut_4_lut (.A(n15016), .B(n15004), .C(\array[201] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3665[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_58_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_58_i6_3_lut_4_lut (.A(n15016), .B(n15004), .C(\array[201] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3665[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_58_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_58_i7_3_lut_4_lut (.A(n15016), .B(n15004), .C(\array[201] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3665[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_58_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_58_i8_3_lut_4_lut (.A(n15016), .B(n15004), .C(\array[201] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3665[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_58_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_57_i1_3_lut_4_lut (.A(n15017), .B(n15004), .C(\array[202] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3673[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_57_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_57_i2_3_lut_4_lut (.A(n15017), .B(n15004), .C(\array[202] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3673[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_57_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_57_i3_3_lut_4_lut (.A(n15017), .B(n15004), .C(\array[202] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3673[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_57_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_57_i4_3_lut_4_lut (.A(n15017), .B(n15004), .C(\array[202] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3673[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_57_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_57_i5_3_lut_4_lut (.A(n15017), .B(n15004), .C(\array[202] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3673[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_57_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_57_i6_3_lut_4_lut (.A(n15017), .B(n15004), .C(\array[202] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3673[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_57_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_57_i7_3_lut_4_lut (.A(n15017), .B(n15004), .C(\array[202] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3673[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_57_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_57_i8_3_lut_4_lut (.A(n15017), .B(n15004), .C(\array[202] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3673[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_57_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_56_i1_3_lut_4_lut (.A(n15018), .B(n15004), .C(\array[203] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3681[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_56_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_56_i2_3_lut_4_lut (.A(n15018), .B(n15004), .C(\array[203] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3681[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_56_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_56_i3_3_lut_4_lut (.A(n15018), .B(n15004), .C(\array[203] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3681[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_56_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_56_i4_3_lut_4_lut (.A(n15018), .B(n15004), .C(\array[203] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3681[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_56_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_56_i5_3_lut_4_lut (.A(n15018), .B(n15004), .C(\array[203] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3681[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_56_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_56_i6_3_lut_4_lut (.A(n15018), .B(n15004), .C(\array[203] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3681[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_56_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_56_i7_3_lut_4_lut (.A(n15018), .B(n15004), .C(\array[203] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3681[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_56_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_56_i8_3_lut_4_lut (.A(n15018), .B(n15004), .C(\array[203] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3681[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_56_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_55_i1_3_lut_4_lut (.A(n15019), .B(n15004), .C(\array[204] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3689[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_55_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_55_i2_3_lut_4_lut (.A(n15019), .B(n15004), .C(\array[204] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3689[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_55_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_55_i3_3_lut_4_lut (.A(n15019), .B(n15004), .C(\array[204] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3689[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_55_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_55_i4_3_lut_4_lut (.A(n15019), .B(n15004), .C(\array[204] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3689[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_55_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_55_i5_3_lut_4_lut (.A(n15019), .B(n15004), .C(\array[204] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3689[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_55_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_55_i6_3_lut_4_lut (.A(n15019), .B(n15004), .C(\array[204] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3689[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_55_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_55_i7_3_lut_4_lut (.A(n15019), .B(n15004), .C(\array[204] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3689[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_55_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_55_i8_3_lut_4_lut (.A(n15019), .B(n15004), .C(\array[204] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3689[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_55_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_54_i1_3_lut_4_lut (.A(n15020), .B(n15004), .C(\array[205] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3697[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_54_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_54_i2_3_lut_4_lut (.A(n15020), .B(n15004), .C(\array[205] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3697[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_54_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_54_i3_3_lut_4_lut (.A(n15020), .B(n15004), .C(\array[205] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3697[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_54_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_54_i4_3_lut_4_lut (.A(n15020), .B(n15004), .C(\array[205] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3697[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_54_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_54_i5_3_lut_4_lut (.A(n15020), .B(n15004), .C(\array[205] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3697[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_54_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_54_i6_3_lut_4_lut (.A(n15020), .B(n15004), .C(\array[205] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3697[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_54_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_54_i7_3_lut_4_lut (.A(n15020), .B(n15004), .C(\array[205] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3697[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_54_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_54_i8_3_lut_4_lut (.A(n15020), .B(n15004), .C(\array[205] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3697[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_54_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_53_i1_3_lut_4_lut (.A(n15021), .B(n15004), .C(\array[206] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3705[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_53_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_53_i2_3_lut_4_lut (.A(n15021), .B(n15004), .C(\array[206] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3705[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_53_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_53_i3_3_lut_4_lut (.A(n15021), .B(n15004), .C(\array[206] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3705[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_53_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_53_i4_3_lut_4_lut (.A(n15021), .B(n15004), .C(\array[206] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3705[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_53_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_53_i5_3_lut_4_lut (.A(n15021), .B(n15004), .C(\array[206] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3705[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_53_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_53_i6_3_lut_4_lut (.A(n15021), .B(n15004), .C(\array[206] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3705[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_53_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_53_i7_3_lut_4_lut (.A(n15021), .B(n15004), .C(\array[206] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3705[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_53_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_53_i8_3_lut_4_lut (.A(n15021), .B(n15004), .C(\array[206] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3705[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_53_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_52_i1_3_lut_4_lut (.A(n15023), .B(n15004), .C(\array[207] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3713[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_52_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_52_i2_3_lut_4_lut (.A(n15023), .B(n15004), .C(\array[207] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3713[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_52_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_52_i3_3_lut_4_lut (.A(n15023), .B(n15004), .C(\array[207] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3713[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_52_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_52_i4_3_lut_4_lut (.A(n15023), .B(n15004), .C(\array[207] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3713[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_52_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_52_i5_3_lut_4_lut (.A(n15023), .B(n15004), .C(\array[207] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3713[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_52_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_52_i6_3_lut_4_lut (.A(n15023), .B(n15004), .C(\array[207] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3713[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_52_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_52_i7_3_lut_4_lut (.A(n15023), .B(n15004), .C(\array[207] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3713[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_52_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_255_i5_3_lut_4_lut (.A(n15011), .B(n14992), .C(\array[4] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2089[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_255_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_52_i8_3_lut_4_lut (.A(n15023), .B(n15004), .C(\array[207] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3713[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_52_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_51_i1_3_lut_4_lut (.A(n15007), .B(n15005), .C(\array[208] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3721[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_51_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i2_3_lut_4_lut (.A(n15007), .B(n15005), .C(\array[208] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3721[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_51_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i3_3_lut_4_lut (.A(n15007), .B(n15005), .C(\array[208] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3721[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_51_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i4_3_lut_4_lut (.A(n15007), .B(n15005), .C(\array[208] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3721[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_51_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i5_3_lut_4_lut (.A(n15007), .B(n15005), .C(\array[208] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3721[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_51_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i6_3_lut_4_lut (.A(n15007), .B(n15005), .C(\array[208] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3721[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_51_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i7_3_lut_4_lut (.A(n15007), .B(n15005), .C(\array[208] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3721[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_51_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_51_i8_3_lut_4_lut (.A(n15007), .B(n15005), .C(\array[208] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3721[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_51_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_50_i1_3_lut_4_lut (.A(n15008), .B(n15005), .C(\array[209] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3729[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_50_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_50_i2_3_lut_4_lut (.A(n15008), .B(n15005), .C(\array[209] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3729[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_50_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_255_i6_3_lut_4_lut (.A(n15011), .B(n14992), .C(\array[4] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2089[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_255_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_50_i3_3_lut_4_lut (.A(n15008), .B(n15005), .C(\array[209] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3729[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_50_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_50_i4_3_lut_4_lut (.A(n15008), .B(n15005), .C(\array[209] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3729[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_50_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_50_i5_3_lut_4_lut (.A(n15008), .B(n15005), .C(\array[209] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3729[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_50_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_50_i6_3_lut_4_lut (.A(n15008), .B(n15005), .C(\array[209] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3729[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_50_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_50_i7_3_lut_4_lut (.A(n15008), .B(n15005), .C(\array[209] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3729[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_50_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_50_i8_3_lut_4_lut (.A(n15008), .B(n15005), .C(\array[209] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3729[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_50_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_49_i1_3_lut_4_lut (.A(n15009), .B(n15005), .C(\array[210] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3737[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_49_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_49_i2_3_lut_4_lut (.A(n15009), .B(n15005), .C(\array[210] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3737[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_49_i2_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i5882 (.BLUT(n14415), .ALUT(n14416), .C0(r_addr[1]), .Z(n14424));
    LUT4 mux_49_i3_3_lut_4_lut (.A(n15009), .B(n15005), .C(\array[210] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3737[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_49_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_49_i4_3_lut_4_lut (.A(n15009), .B(n15005), .C(\array[210] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3737[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_49_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_49_i5_3_lut_4_lut (.A(n15009), .B(n15005), .C(\array[210] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3737[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_49_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_49_i6_3_lut_4_lut (.A(n15009), .B(n15005), .C(\array[210] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3737[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_49_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_49_i7_3_lut_4_lut (.A(n15009), .B(n15005), .C(\array[210] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3737[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_49_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_49_i8_3_lut_4_lut (.A(n15009), .B(n15005), .C(\array[210] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3737[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_49_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_48_i1_3_lut_4_lut (.A(n15010), .B(n15005), .C(\array[211] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3745[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_48_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_48_i2_3_lut_4_lut (.A(n15010), .B(n15005), .C(\array[211] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3745[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_48_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_48_i3_3_lut_4_lut (.A(n15010), .B(n15005), .C(\array[211] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3745[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_48_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_48_i4_3_lut_4_lut (.A(n15010), .B(n15005), .C(\array[211] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3745[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_48_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_48_i5_3_lut_4_lut (.A(n15010), .B(n15005), .C(\array[211] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3745[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_48_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_48_i6_3_lut_4_lut (.A(n15010), .B(n15005), .C(\array[211] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3745[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_48_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_48_i7_3_lut_4_lut (.A(n15010), .B(n15005), .C(\array[211] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3745[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_48_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_48_i8_3_lut_4_lut (.A(n15010), .B(n15005), .C(\array[211] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3745[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_48_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_47_i1_3_lut_4_lut (.A(n15011), .B(n15005), .C(\array[212] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3753[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_47_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_47_i2_3_lut_4_lut (.A(n15011), .B(n15005), .C(\array[212] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3753[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_47_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_47_i3_3_lut_4_lut (.A(n15011), .B(n15005), .C(\array[212] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3753[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_47_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_47_i4_3_lut_4_lut (.A(n15011), .B(n15005), .C(\array[212] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3753[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_47_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_47_i5_3_lut_4_lut (.A(n15011), .B(n15005), .C(\array[212] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3753[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_47_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_47_i6_3_lut_4_lut (.A(n15011), .B(n15005), .C(\array[212] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3753[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_47_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_47_i7_3_lut_4_lut (.A(n15011), .B(n15005), .C(\array[212] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3753[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_47_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_47_i8_3_lut_4_lut (.A(n15011), .B(n15005), .C(\array[212] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3753[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_47_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_46_i1_3_lut_4_lut (.A(n15012), .B(n15005), .C(\array[213] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3761[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_46_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_46_i2_3_lut_4_lut (.A(n15012), .B(n15005), .C(\array[213] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3761[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_46_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_46_i3_3_lut_4_lut (.A(n15012), .B(n15005), .C(\array[213] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3761[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_46_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_46_i4_3_lut_4_lut (.A(n15012), .B(n15005), .C(\array[213] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3761[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_46_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_46_i5_3_lut_4_lut (.A(n15012), .B(n15005), .C(\array[213] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3761[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_46_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_46_i6_3_lut_4_lut (.A(n15012), .B(n15005), .C(\array[213] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3761[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_46_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_46_i7_3_lut_4_lut (.A(n15012), .B(n15005), .C(\array[213] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3761[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_46_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_46_i8_3_lut_4_lut (.A(n15012), .B(n15005), .C(\array[213] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3761[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_46_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_45_i1_3_lut_4_lut (.A(n15013), .B(n15005), .C(\array[214] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3769[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_45_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_255_i7_3_lut_4_lut (.A(n15011), .B(n14992), .C(\array[4] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2089[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_255_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_45_i2_3_lut_4_lut (.A(n15013), .B(n15005), .C(\array[214] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3769[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_45_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_45_i3_3_lut_4_lut (.A(n15013), .B(n15005), .C(\array[214] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3769[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_45_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_45_i4_3_lut_4_lut (.A(n15013), .B(n15005), .C(\array[214] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3769[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_45_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_45_i5_3_lut_4_lut (.A(n15013), .B(n15005), .C(\array[214] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3769[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_45_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_45_i6_3_lut_4_lut (.A(n15013), .B(n15005), .C(\array[214] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3769[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_45_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_45_i7_3_lut_4_lut (.A(n15013), .B(n15005), .C(\array[214] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3769[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_45_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_45_i8_3_lut_4_lut (.A(n15013), .B(n15005), .C(\array[214] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3769[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_45_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_44_i1_3_lut_4_lut (.A(n15014), .B(n15005), .C(\array[215] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3777[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_44_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_44_i2_3_lut_4_lut (.A(n15014), .B(n15005), .C(\array[215] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3777[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_44_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_44_i3_3_lut_4_lut (.A(n15014), .B(n15005), .C(\array[215] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3777[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_44_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_44_i4_3_lut_4_lut (.A(n15014), .B(n15005), .C(\array[215] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3777[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_44_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_44_i5_3_lut_4_lut (.A(n15014), .B(n15005), .C(\array[215] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3777[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_44_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_44_i6_3_lut_4_lut (.A(n15014), .B(n15005), .C(\array[215] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3777[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_44_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_44_i7_3_lut_4_lut (.A(n15014), .B(n15005), .C(\array[215] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3777[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_44_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_44_i8_3_lut_4_lut (.A(n15014), .B(n15005), .C(\array[215] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3777[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_44_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_43_i1_3_lut_4_lut (.A(n15015), .B(n15005), .C(\array[216] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3785[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_43_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_43_i2_3_lut_4_lut (.A(n15015), .B(n15005), .C(\array[216] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3785[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_43_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_43_i3_3_lut_4_lut (.A(n15015), .B(n15005), .C(\array[216] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3785[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_43_i3_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i5341 (.BLUT(n13874), .ALUT(n13875), .C0(r_addr[1]), .Z(n13883));
    LUT4 mux_43_i4_3_lut_4_lut (.A(n15015), .B(n15005), .C(\array[216] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3785[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_43_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_43_i5_3_lut_4_lut (.A(n15015), .B(n15005), .C(\array[216] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3785[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_43_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_43_i6_3_lut_4_lut (.A(n15015), .B(n15005), .C(\array[216] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3785[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_43_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_43_i7_3_lut_4_lut (.A(n15015), .B(n15005), .C(\array[216] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3785[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_43_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_43_i8_3_lut_4_lut (.A(n15015), .B(n15005), .C(\array[216] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3785[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_43_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_42_i1_3_lut_4_lut (.A(n15016), .B(n15005), .C(\array[217] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3793[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_42_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_42_i2_3_lut_4_lut (.A(n15016), .B(n15005), .C(\array[217] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3793[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_42_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_42_i3_3_lut_4_lut (.A(n15016), .B(n15005), .C(\array[217] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3793[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_42_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_42_i4_3_lut_4_lut (.A(n15016), .B(n15005), .C(\array[217] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3793[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_42_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_42_i5_3_lut_4_lut (.A(n15016), .B(n15005), .C(\array[217] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3793[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_42_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_42_i6_3_lut_4_lut (.A(n15016), .B(n15005), .C(\array[217] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3793[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_42_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_42_i7_3_lut_4_lut (.A(n15016), .B(n15005), .C(\array[217] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3793[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_42_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_42_i8_3_lut_4_lut (.A(n15016), .B(n15005), .C(\array[217] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3793[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_42_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_41_i1_3_lut_4_lut (.A(n15017), .B(n15005), .C(\array[218] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3801[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_41_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_41_i2_3_lut_4_lut (.A(n15017), .B(n15005), .C(\array[218] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3801[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_41_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_41_i3_3_lut_4_lut (.A(n15017), .B(n15005), .C(\array[218] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3801[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_41_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_41_i4_3_lut_4_lut (.A(n15017), .B(n15005), .C(\array[218] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3801[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_41_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_41_i5_3_lut_4_lut (.A(n15017), .B(n15005), .C(\array[218] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3801[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_41_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_41_i6_3_lut_4_lut (.A(n15017), .B(n15005), .C(\array[218] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3801[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_41_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_41_i7_3_lut_4_lut (.A(n15017), .B(n15005), .C(\array[218] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3801[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_41_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_41_i8_3_lut_4_lut (.A(n15017), .B(n15005), .C(\array[218] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3801[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_41_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_40_i1_3_lut_4_lut (.A(n15018), .B(n15005), .C(\array[219] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3809[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_40_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_40_i2_3_lut_4_lut (.A(n15018), .B(n15005), .C(\array[219] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3809[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_40_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_40_i3_3_lut_4_lut (.A(n15018), .B(n15005), .C(\array[219] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3809[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_40_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_40_i4_3_lut_4_lut (.A(n15018), .B(n15005), .C(\array[219] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3809[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_40_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_40_i5_3_lut_4_lut (.A(n15018), .B(n15005), .C(\array[219] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3809[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_40_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_40_i6_3_lut_4_lut (.A(n15018), .B(n15005), .C(\array[219] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3809[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_40_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_40_i7_3_lut_4_lut (.A(n15018), .B(n15005), .C(\array[219] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3809[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_40_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_40_i8_3_lut_4_lut (.A(n15018), .B(n15005), .C(\array[219] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3809[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_40_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_39_i1_3_lut_4_lut (.A(n15019), .B(n15005), .C(\array[220] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3817[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_39_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_39_i2_3_lut_4_lut (.A(n15019), .B(n15005), .C(\array[220] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3817[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_39_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_39_i3_3_lut_4_lut (.A(n15019), .B(n15005), .C(\array[220] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3817[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_39_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_39_i4_3_lut_4_lut (.A(n15019), .B(n15005), .C(\array[220] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3817[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_39_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_39_i5_3_lut_4_lut (.A(n15019), .B(n15005), .C(\array[220] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3817[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_39_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_39_i6_3_lut_4_lut (.A(n15019), .B(n15005), .C(\array[220] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3817[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_39_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_39_i7_3_lut_4_lut (.A(n15019), .B(n15005), .C(\array[220] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3817[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_39_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_39_i8_3_lut_4_lut (.A(n15019), .B(n15005), .C(\array[220] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3817[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_39_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_38_i1_3_lut_4_lut (.A(n15020), .B(n15005), .C(\array[221] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3825[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_38_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_38_i2_3_lut_4_lut (.A(n15020), .B(n15005), .C(\array[221] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3825[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_38_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_38_i3_3_lut_4_lut (.A(n15020), .B(n15005), .C(\array[221] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3825[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_38_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_38_i4_3_lut_4_lut (.A(n15020), .B(n15005), .C(\array[221] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3825[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_38_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_38_i5_3_lut_4_lut (.A(n15020), .B(n15005), .C(\array[221] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3825[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_38_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_38_i6_3_lut_4_lut (.A(n15020), .B(n15005), .C(\array[221] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3825[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_38_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_38_i7_3_lut_4_lut (.A(n15020), .B(n15005), .C(\array[221] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3825[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_38_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_38_i8_3_lut_4_lut (.A(n15020), .B(n15005), .C(\array[221] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3825[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_38_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_37_i1_3_lut_4_lut (.A(n15021), .B(n15005), .C(\array[222] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3833[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_37_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_37_i2_3_lut_4_lut (.A(n15021), .B(n15005), .C(\array[222] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3833[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_37_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_37_i3_3_lut_4_lut (.A(n15021), .B(n15005), .C(\array[222] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3833[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_37_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_37_i4_3_lut_4_lut (.A(n15021), .B(n15005), .C(\array[222] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3833[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_37_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_37_i5_3_lut_4_lut (.A(n15021), .B(n15005), .C(\array[222] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3833[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_37_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_37_i6_3_lut_4_lut (.A(n15021), .B(n15005), .C(\array[222] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3833[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_37_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_37_i7_3_lut_4_lut (.A(n15021), .B(n15005), .C(\array[222] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3833[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_37_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_37_i8_3_lut_4_lut (.A(n15021), .B(n15005), .C(\array[222] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3833[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_37_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_36_i1_3_lut_4_lut (.A(n15023), .B(n15005), .C(\array[223] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3841[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_36_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_36_i2_3_lut_4_lut (.A(n15023), .B(n15005), .C(\array[223] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3841[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_36_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_255_i8_3_lut_4_lut (.A(n15011), .B(n14992), .C(\array[4] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2089[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_255_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_36_i3_3_lut_4_lut (.A(n15023), .B(n15005), .C(\array[223] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3841[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_36_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_36_i4_3_lut_4_lut (.A(n15023), .B(n15005), .C(\array[223] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3841[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_36_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_36_i5_3_lut_4_lut (.A(n15023), .B(n15005), .C(\array[223] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3841[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_36_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_36_i6_3_lut_4_lut (.A(n15023), .B(n15005), .C(\array[223] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3841[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_36_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_36_i7_3_lut_4_lut (.A(n15023), .B(n15005), .C(\array[223] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3841[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_36_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_36_i8_3_lut_4_lut (.A(n15023), .B(n15005), .C(\array[223] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3841[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_36_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_35_i1_3_lut_4_lut (.A(n15007), .B(n15006), .C(\array[224] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3849[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_35_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_35_i2_3_lut_4_lut (.A(n15007), .B(n15006), .C(\array[224] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3849[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_35_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_35_i3_3_lut_4_lut (.A(n15007), .B(n15006), .C(\array[224] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3849[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_35_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_35_i4_3_lut_4_lut (.A(n15007), .B(n15006), .C(\array[224] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3849[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_35_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_35_i5_3_lut_4_lut (.A(n15007), .B(n15006), .C(\array[224] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3849[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_35_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_35_i6_3_lut_4_lut (.A(n15007), .B(n15006), .C(\array[224] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3849[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_35_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_35_i7_3_lut_4_lut (.A(n15007), .B(n15006), .C(\array[224] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3849[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_35_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_35_i8_3_lut_4_lut (.A(n15007), .B(n15006), .C(\array[224] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3849[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_35_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_34_i1_3_lut_4_lut (.A(n15008), .B(n15006), .C(\array[225] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3857[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_34_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_34_i2_3_lut_4_lut (.A(n15008), .B(n15006), .C(\array[225] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3857[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_34_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_34_i3_3_lut_4_lut (.A(n15008), .B(n15006), .C(\array[225] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3857[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_34_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_34_i4_3_lut_4_lut (.A(n15008), .B(n15006), .C(\array[225] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3857[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_34_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_34_i5_3_lut_4_lut (.A(n15008), .B(n15006), .C(\array[225] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3857[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_34_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_34_i6_3_lut_4_lut (.A(n15008), .B(n15006), .C(\array[225] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3857[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_34_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_34_i7_3_lut_4_lut (.A(n15008), .B(n15006), .C(\array[225] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3857[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_34_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_34_i8_3_lut_4_lut (.A(n15008), .B(n15006), .C(\array[225] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3857[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_34_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_33_i1_3_lut_4_lut (.A(n15009), .B(n15006), .C(\array[226] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3865[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_33_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_33_i2_3_lut_4_lut (.A(n15009), .B(n15006), .C(\array[226] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3865[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_33_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_33_i3_3_lut_4_lut (.A(n15009), .B(n15006), .C(\array[226] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3865[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_33_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_33_i4_3_lut_4_lut (.A(n15009), .B(n15006), .C(\array[226] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3865[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_33_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_33_i5_3_lut_4_lut (.A(n15009), .B(n15006), .C(\array[226] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3865[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_33_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_33_i6_3_lut_4_lut (.A(n15009), .B(n15006), .C(\array[226] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3865[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_33_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_33_i7_3_lut_4_lut (.A(n15009), .B(n15006), .C(\array[226] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3865[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_33_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_33_i8_3_lut_4_lut (.A(n15009), .B(n15006), .C(\array[226] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3865[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_33_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_32_i1_3_lut_4_lut (.A(n15010), .B(n15006), .C(\array[227] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3873[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_32_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_32_i2_3_lut_4_lut (.A(n15010), .B(n15006), .C(\array[227] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3873[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_32_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_32_i3_3_lut_4_lut (.A(n15010), .B(n15006), .C(\array[227] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3873[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_32_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_32_i4_3_lut_4_lut (.A(n15010), .B(n15006), .C(\array[227] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3873[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_32_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_32_i5_3_lut_4_lut (.A(n15010), .B(n15006), .C(\array[227] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3873[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_32_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_32_i6_3_lut_4_lut (.A(n15010), .B(n15006), .C(\array[227] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3873[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_32_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_32_i7_3_lut_4_lut (.A(n15010), .B(n15006), .C(\array[227] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3873[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_32_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_32_i8_3_lut_4_lut (.A(n15010), .B(n15006), .C(\array[227] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3873[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_32_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_31_i1_3_lut_4_lut (.A(n15011), .B(n15006), .C(\array[228] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3881[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_31_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_31_i2_3_lut_4_lut (.A(n15011), .B(n15006), .C(\array[228] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3881[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_31_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_31_i3_3_lut_4_lut (.A(n15011), .B(n15006), .C(\array[228] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3881[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_31_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_31_i4_3_lut_4_lut (.A(n15011), .B(n15006), .C(\array[228] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3881[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_31_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_31_i5_3_lut_4_lut (.A(n15011), .B(n15006), .C(\array[228] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3881[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_31_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_31_i6_3_lut_4_lut (.A(n15011), .B(n15006), .C(\array[228] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3881[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_31_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_31_i7_3_lut_4_lut (.A(n15011), .B(n15006), .C(\array[228] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3881[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_31_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_31_i8_3_lut_4_lut (.A(n15011), .B(n15006), .C(\array[228] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3881[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_31_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_30_i1_3_lut_4_lut (.A(n15012), .B(n15006), .C(\array[229] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3889[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_30_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_30_i2_3_lut_4_lut (.A(n15012), .B(n15006), .C(\array[229] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3889[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_30_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_30_i3_3_lut_4_lut (.A(n15012), .B(n15006), .C(\array[229] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3889[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_30_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_30_i4_3_lut_4_lut (.A(n15012), .B(n15006), .C(\array[229] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3889[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_30_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_30_i5_3_lut_4_lut (.A(n15012), .B(n15006), .C(\array[229] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3889[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_30_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_30_i6_3_lut_4_lut (.A(n15012), .B(n15006), .C(\array[229] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3889[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_30_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_30_i7_3_lut_4_lut (.A(n15012), .B(n15006), .C(\array[229] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3889[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_30_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_30_i8_3_lut_4_lut (.A(n15012), .B(n15006), .C(\array[229] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3889[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_30_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_29_i1_3_lut_4_lut (.A(n15013), .B(n15006), .C(\array[230] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3897[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_29_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_29_i2_3_lut_4_lut (.A(n15013), .B(n15006), .C(\array[230] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3897[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_29_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_29_i3_3_lut_4_lut (.A(n15013), .B(n15006), .C(\array[230] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3897[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_29_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_29_i4_3_lut_4_lut (.A(n15013), .B(n15006), .C(\array[230] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3897[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_29_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_29_i5_3_lut_4_lut (.A(n15013), .B(n15006), .C(\array[230] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3897[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_29_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_29_i6_3_lut_4_lut (.A(n15013), .B(n15006), .C(\array[230] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3897[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_29_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_29_i7_3_lut_4_lut (.A(n15013), .B(n15006), .C(\array[230] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3897[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_29_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_29_i8_3_lut_4_lut (.A(n15013), .B(n15006), .C(\array[230] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3897[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_29_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_28_i1_3_lut_4_lut (.A(n15014), .B(n15006), .C(\array[231] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3905[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_28_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_28_i2_3_lut_4_lut (.A(n15014), .B(n15006), .C(\array[231] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3905[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_28_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_28_i3_3_lut_4_lut (.A(n15014), .B(n15006), .C(\array[231] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3905[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_28_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_28_i4_3_lut_4_lut (.A(n15014), .B(n15006), .C(\array[231] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3905[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_28_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_28_i5_3_lut_4_lut (.A(n15014), .B(n15006), .C(\array[231] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3905[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_28_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_28_i6_3_lut_4_lut (.A(n15014), .B(n15006), .C(\array[231] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3905[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_28_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_254_i1_3_lut_4_lut (.A(n15012), .B(n14992), .C(\array[5] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2097[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_254_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_28_i7_3_lut_4_lut (.A(n15014), .B(n15006), .C(\array[231] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3905[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_28_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_28_i8_3_lut_4_lut (.A(n15014), .B(n15006), .C(\array[231] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3905[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_28_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_27_i1_3_lut_4_lut (.A(n15015), .B(n15006), .C(\array[232] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3913[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_27_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_27_i2_3_lut_4_lut (.A(n15015), .B(n15006), .C(\array[232] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3913[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_27_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_27_i3_3_lut_4_lut (.A(n15015), .B(n15006), .C(\array[232] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3913[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_27_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_27_i4_3_lut_4_lut (.A(n15015), .B(n15006), .C(\array[232] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3913[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_27_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_27_i5_3_lut_4_lut (.A(n15015), .B(n15006), .C(\array[232] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3913[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_27_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_27_i6_3_lut_4_lut (.A(n15015), .B(n15006), .C(\array[232] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3913[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_27_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_27_i7_3_lut_4_lut (.A(n15015), .B(n15006), .C(\array[232] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3913[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_27_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_27_i8_3_lut_4_lut (.A(n15015), .B(n15006), .C(\array[232] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3913[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_27_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_26_i1_3_lut_4_lut (.A(n15016), .B(n15006), .C(\array[233] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3921[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_26_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_26_i2_3_lut_4_lut (.A(n15016), .B(n15006), .C(\array[233] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3921[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_26_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_26_i3_3_lut_4_lut (.A(n15016), .B(n15006), .C(\array[233] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3921[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_26_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_26_i4_3_lut_4_lut (.A(n15016), .B(n15006), .C(\array[233] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3921[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_26_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_26_i5_3_lut_4_lut (.A(n15016), .B(n15006), .C(\array[233] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3921[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_26_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_26_i6_3_lut_4_lut (.A(n15016), .B(n15006), .C(\array[233] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3921[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_26_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_26_i7_3_lut_4_lut (.A(n15016), .B(n15006), .C(\array[233] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3921[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_26_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_26_i8_3_lut_4_lut (.A(n15016), .B(n15006), .C(\array[233] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3921[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_26_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_25_i1_3_lut_4_lut (.A(n15017), .B(n15006), .C(\array[234] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3929[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_25_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_25_i2_3_lut_4_lut (.A(n15017), .B(n15006), .C(\array[234] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3929[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_25_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_25_i3_3_lut_4_lut (.A(n15017), .B(n15006), .C(\array[234] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3929[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_25_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_25_i4_3_lut_4_lut (.A(n15017), .B(n15006), .C(\array[234] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3929[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_25_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_25_i5_3_lut_4_lut (.A(n15017), .B(n15006), .C(\array[234] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3929[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_25_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_25_i6_3_lut_4_lut (.A(n15017), .B(n15006), .C(\array[234] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3929[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_25_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_25_i7_3_lut_4_lut (.A(n15017), .B(n15006), .C(\array[234] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3929[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_25_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_25_i8_3_lut_4_lut (.A(n15017), .B(n15006), .C(\array[234] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3929[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_25_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_24_i1_3_lut_4_lut (.A(n15018), .B(n15006), .C(\array[235] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3937[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_24_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_24_i2_3_lut_4_lut (.A(n15018), .B(n15006), .C(\array[235] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3937[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_24_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_24_i3_3_lut_4_lut (.A(n15018), .B(n15006), .C(\array[235] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3937[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_24_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_24_i4_3_lut_4_lut (.A(n15018), .B(n15006), .C(\array[235] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3937[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_24_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_24_i5_3_lut_4_lut (.A(n15018), .B(n15006), .C(\array[235] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3937[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_24_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_24_i6_3_lut_4_lut (.A(n15018), .B(n15006), .C(\array[235] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3937[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_24_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_254_i2_3_lut_4_lut (.A(n15012), .B(n14992), .C(\array[5] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2097[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_254_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_24_i7_3_lut_4_lut (.A(n15018), .B(n15006), .C(\array[235] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3937[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_24_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_24_i8_3_lut_4_lut (.A(n15018), .B(n15006), .C(\array[235] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3937[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_24_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i1_3_lut_4_lut (.A(n15019), .B(n15006), .C(\array[236] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3945[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_23_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i2_3_lut_4_lut (.A(n15019), .B(n15006), .C(\array[236] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3945[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_23_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i3_3_lut_4_lut (.A(n15019), .B(n15006), .C(\array[236] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3945[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_23_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_254_i3_3_lut_4_lut (.A(n15012), .B(n14992), .C(\array[5] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2097[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_254_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i4_3_lut_4_lut (.A(n15019), .B(n15006), .C(\array[236] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3945[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_23_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_254_i4_3_lut_4_lut (.A(n15012), .B(n14992), .C(\array[5] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2097[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_254_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i5_3_lut_4_lut (.A(n15019), .B(n15006), .C(\array[236] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3945[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_23_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i6_3_lut_4_lut (.A(n15019), .B(n15006), .C(\array[236] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3945[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_23_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i7_3_lut_4_lut (.A(n15019), .B(n15006), .C(\array[236] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3945[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_23_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_23_i8_3_lut_4_lut (.A(n15019), .B(n15006), .C(\array[236] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3945[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_23_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i1_3_lut_4_lut (.A(n15020), .B(n15006), .C(\array[237] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3953[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_22_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i2_3_lut_4_lut (.A(n15020), .B(n15006), .C(\array[237] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3953[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_22_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i3_3_lut_4_lut (.A(n15020), .B(n15006), .C(\array[237] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3953[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_22_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_254_i5_3_lut_4_lut (.A(n15012), .B(n14992), .C(\array[5] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2097[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_254_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_254_i6_3_lut_4_lut (.A(n15012), .B(n14992), .C(\array[5] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2097[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_254_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i4_3_lut_4_lut (.A(n15020), .B(n15006), .C(\array[237] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3953[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_22_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i5_3_lut_4_lut (.A(n15020), .B(n15006), .C(\array[237] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3953[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_22_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_254_i7_3_lut_4_lut (.A(n15012), .B(n14992), .C(\array[5] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2097[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_254_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i6_3_lut_4_lut (.A(n15020), .B(n15006), .C(\array[237] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3953[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_22_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_254_i8_3_lut_4_lut (.A(n15012), .B(n14992), .C(\array[5] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2097[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_254_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i7_3_lut_4_lut (.A(n15020), .B(n15006), .C(\array[237] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3953[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_22_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_22_i8_3_lut_4_lut (.A(n15020), .B(n15006), .C(\array[237] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3953[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_22_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i1_3_lut_4_lut (.A(n15021), .B(n15006), .C(\array[238] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3961[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_21_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i2_3_lut_4_lut (.A(n15021), .B(n15006), .C(\array[238] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3961[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_21_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i3_3_lut_4_lut (.A(n15021), .B(n15006), .C(\array[238] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3961[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_21_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i4_3_lut_4_lut (.A(n15021), .B(n15006), .C(\array[238] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3961[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_21_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i5_3_lut_4_lut (.A(n15021), .B(n15006), .C(\array[238] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3961[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_21_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i6_3_lut_4_lut (.A(n15021), .B(n15006), .C(\array[238] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3961[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_21_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_253_i1_3_lut_4_lut (.A(n15013), .B(n14992), .C(\array[6] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2105[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_253_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i7_3_lut_4_lut (.A(n15021), .B(n15006), .C(\array[238] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3961[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_21_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_21_i8_3_lut_4_lut (.A(n15021), .B(n15006), .C(\array[238] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3961[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_21_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_20_i1_3_lut_4_lut (.A(n15023), .B(n15006), .C(\array[239] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3969[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_20_i1_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i2_3_lut_4_lut (.A(n15023), .B(n15006), .C(\array[239] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3969[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_20_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i3_3_lut_4_lut (.A(n15023), .B(n15006), .C(\array[239] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3969[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_20_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i4_3_lut_4_lut (.A(n15023), .B(n15006), .C(\array[239] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3969[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_20_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i5_3_lut_4_lut (.A(n15023), .B(n15006), .C(\array[239] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3969[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_20_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i6_3_lut_4_lut (.A(n15023), .B(n15006), .C(\array[239] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3969[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_20_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i7_3_lut_4_lut (.A(n15023), .B(n15006), .C(\array[239] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3969[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_20_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_20_i8_3_lut_4_lut (.A(n15023), .B(n15006), .C(\array[239] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3969[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_20_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_19_i1_3_lut_4_lut (.A(n15007), .B(n15022), .C(\array[240] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3977[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_19_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_19_i2_3_lut_4_lut (.A(n15007), .B(n15022), .C(\array[240] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3977[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_19_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_19_i3_3_lut_4_lut (.A(n15007), .B(n15022), .C(\array[240] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3977[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_19_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_19_i4_3_lut_4_lut (.A(n15007), .B(n15022), .C(\array[240] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3977[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_19_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_19_i5_3_lut_4_lut (.A(n15007), .B(n15022), .C(\array[240] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3977[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_19_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_19_i6_3_lut_4_lut (.A(n15007), .B(n15022), .C(\array[240] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3977[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_19_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_19_i7_3_lut_4_lut (.A(n15007), .B(n15022), .C(\array[240] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3977[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_19_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_19_i8_3_lut_4_lut (.A(n15007), .B(n15022), .C(\array[240] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3977[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_19_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_18_i1_3_lut_4_lut (.A(n15008), .B(n15022), .C(\array[241] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3985[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_18_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_18_i2_3_lut_4_lut (.A(n15008), .B(n15022), .C(\array[241] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3985[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_18_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_18_i3_3_lut_4_lut (.A(n15008), .B(n15022), .C(\array[241] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3985[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_18_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_18_i4_3_lut_4_lut (.A(n15008), .B(n15022), .C(\array[241] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3985[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_18_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_18_i5_3_lut_4_lut (.A(n15008), .B(n15022), .C(\array[241] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3985[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_18_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_18_i6_3_lut_4_lut (.A(n15008), .B(n15022), .C(\array[241] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3985[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_18_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_18_i7_3_lut_4_lut (.A(n15008), .B(n15022), .C(\array[241] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3985[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_18_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_18_i8_3_lut_4_lut (.A(n15008), .B(n15022), .C(\array[241] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3985[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_18_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_17_i1_3_lut_4_lut (.A(n15009), .B(n15022), .C(\array[242] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_3993[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_17_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_17_i2_3_lut_4_lut (.A(n15009), .B(n15022), .C(\array[242] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_3993[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_17_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_17_i3_3_lut_4_lut (.A(n15009), .B(n15022), .C(\array[242] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_3993[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_17_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_17_i4_3_lut_4_lut (.A(n15009), .B(n15022), .C(\array[242] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_3993[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_17_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_17_i5_3_lut_4_lut (.A(n15009), .B(n15022), .C(\array[242] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_3993[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_17_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_17_i6_3_lut_4_lut (.A(n15009), .B(n15022), .C(\array[242] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_3993[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_17_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_17_i7_3_lut_4_lut (.A(n15009), .B(n15022), .C(\array[242] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_3993[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_17_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_17_i8_3_lut_4_lut (.A(n15009), .B(n15022), .C(\array[242] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_3993[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_17_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_16_i1_3_lut_4_lut (.A(n15010), .B(n15022), .C(\array[243] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_4001[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_16_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_16_i2_3_lut_4_lut (.A(n15010), .B(n15022), .C(\array[243] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_4001[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_16_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_16_i3_3_lut_4_lut (.A(n15010), .B(n15022), .C(\array[243] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_4001[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_16_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_16_i4_3_lut_4_lut (.A(n15010), .B(n15022), .C(\array[243] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_4001[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_16_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_16_i5_3_lut_4_lut (.A(n15010), .B(n15022), .C(\array[243] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_4001[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_16_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_16_i6_3_lut_4_lut (.A(n15010), .B(n15022), .C(\array[243] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_4001[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_16_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_16_i7_3_lut_4_lut (.A(n15010), .B(n15022), .C(\array[243] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_4001[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_16_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_16_i8_3_lut_4_lut (.A(n15010), .B(n15022), .C(\array[243] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_4001[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_16_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_15_i1_3_lut_4_lut (.A(n15011), .B(n15022), .C(\array[244] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_4009[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_15_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_15_i2_3_lut_4_lut (.A(n15011), .B(n15022), .C(\array[244] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_4009[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_15_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_15_i3_3_lut_4_lut (.A(n15011), .B(n15022), .C(\array[244] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_4009[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_15_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_15_i4_3_lut_4_lut (.A(n15011), .B(n15022), .C(\array[244] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_4009[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_15_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_15_i5_3_lut_4_lut (.A(n15011), .B(n15022), .C(\array[244] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_4009[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_15_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_15_i6_3_lut_4_lut (.A(n15011), .B(n15022), .C(\array[244] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_4009[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_15_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_15_i7_3_lut_4_lut (.A(n15011), .B(n15022), .C(\array[244] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_4009[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_15_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_15_i8_3_lut_4_lut (.A(n15011), .B(n15022), .C(\array[244] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_4009[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_15_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_14_i1_3_lut_4_lut (.A(n15012), .B(n15022), .C(\array[245] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_4017[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_14_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_14_i2_3_lut_4_lut (.A(n15012), .B(n15022), .C(\array[245] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_4017[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_14_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_14_i3_3_lut_4_lut (.A(n15012), .B(n15022), .C(\array[245] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_4017[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_14_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_14_i4_3_lut_4_lut (.A(n15012), .B(n15022), .C(\array[245] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_4017[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_14_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_14_i5_3_lut_4_lut (.A(n15012), .B(n15022), .C(\array[245] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_4017[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_14_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_14_i6_3_lut_4_lut (.A(n15012), .B(n15022), .C(\array[245] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_4017[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_14_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_14_i7_3_lut_4_lut (.A(n15012), .B(n15022), .C(\array[245] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_4017[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_14_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_14_i8_3_lut_4_lut (.A(n15012), .B(n15022), .C(\array[245] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_4017[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_14_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_13_i1_3_lut_4_lut (.A(n15013), .B(n15022), .C(\array[246] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_4025[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_13_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_13_i2_3_lut_4_lut (.A(n15013), .B(n15022), .C(\array[246] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_4025[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_13_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_13_i3_3_lut_4_lut (.A(n15013), .B(n15022), .C(\array[246] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_4025[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_13_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_13_i4_3_lut_4_lut (.A(n15013), .B(n15022), .C(\array[246] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_4025[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_13_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_13_i5_3_lut_4_lut (.A(n15013), .B(n15022), .C(\array[246] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_4025[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_13_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_13_i6_3_lut_4_lut (.A(n15013), .B(n15022), .C(\array[246] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_4025[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_13_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_13_i7_3_lut_4_lut (.A(n15013), .B(n15022), .C(\array[246] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_4025[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_13_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_13_i8_3_lut_4_lut (.A(n15013), .B(n15022), .C(\array[246] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_4025[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_13_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_12_i1_3_lut_4_lut (.A(n15014), .B(n15022), .C(\array[247] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_4033[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_12_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_12_i2_3_lut_4_lut (.A(n15014), .B(n15022), .C(\array[247] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_4033[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_12_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_12_i3_3_lut_4_lut (.A(n15014), .B(n15022), .C(\array[247] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_4033[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_12_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_12_i4_3_lut_4_lut (.A(n15014), .B(n15022), .C(\array[247] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_4033[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_12_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_12_i5_3_lut_4_lut (.A(n15014), .B(n15022), .C(\array[247] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_4033[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_12_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_12_i6_3_lut_4_lut (.A(n15014), .B(n15022), .C(\array[247] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_4033[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_12_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_12_i7_3_lut_4_lut (.A(n15014), .B(n15022), .C(\array[247] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_4033[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_12_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_12_i8_3_lut_4_lut (.A(n15014), .B(n15022), .C(\array[247] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_4033[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_12_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i1_3_lut_4_lut (.A(n15015), .B(n15022), .C(\array[248] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_4041[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_11_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i2_3_lut_4_lut (.A(n15015), .B(n15022), .C(\array[248] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_4041[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_11_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i3_3_lut_4_lut (.A(n15015), .B(n15022), .C(\array[248] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_4041[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_11_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i4_3_lut_4_lut (.A(n15015), .B(n15022), .C(\array[248] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_4041[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_11_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i5_3_lut_4_lut (.A(n15015), .B(n15022), .C(\array[248] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_4041[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_11_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i6_3_lut_4_lut (.A(n15015), .B(n15022), .C(\array[248] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_4041[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_11_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i7_3_lut_4_lut (.A(n15015), .B(n15022), .C(\array[248] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_4041[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_11_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_11_i8_3_lut_4_lut (.A(n15015), .B(n15022), .C(\array[248] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_4041[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_11_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i1_3_lut_4_lut (.A(n15016), .B(n15022), .C(\array[249] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_4049[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_10_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i2_3_lut_4_lut (.A(n15016), .B(n15022), .C(\array[249] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_4049[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_10_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i3_3_lut_4_lut (.A(n15016), .B(n15022), .C(\array[249] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_4049[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_10_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i4_3_lut_4_lut (.A(n15016), .B(n15022), .C(\array[249] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_4049[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_10_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i5_3_lut_4_lut (.A(n15016), .B(n15022), .C(\array[249] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_4049[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_10_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i6_3_lut_4_lut (.A(n15016), .B(n15022), .C(\array[249] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_4049[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_10_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i7_3_lut_4_lut (.A(n15016), .B(n15022), .C(\array[249] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_4049[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_10_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_10_i8_3_lut_4_lut (.A(n15016), .B(n15022), .C(\array[249] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_4049[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_10_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i1_3_lut_4_lut (.A(n15017), .B(n15022), .C(\array[250] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_4057[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i2_3_lut_4_lut (.A(n15017), .B(n15022), .C(\array[250] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_4057[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i3_3_lut_4_lut (.A(n15017), .B(n15022), .C(\array[250] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_4057[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n15017), .B(n15022), .C(\array[250] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_4057[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i5_3_lut_4_lut (.A(n15017), .B(n15022), .C(\array[250] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_4057[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n15017), .B(n15022), .C(\array[250] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_4057[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n15017), .B(n15022), .C(\array[250] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_4057[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n15017), .B(n15022), .C(\array[250] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_4057[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_8_i1_3_lut_4_lut (.A(n15018), .B(n15022), .C(\array[251] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_4065[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_8_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_8_i2_3_lut_4_lut (.A(n15018), .B(n15022), .C(\array[251] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_4065[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_8_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_8_i3_3_lut_4_lut (.A(n15018), .B(n15022), .C(\array[251] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_4065[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_8_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_8_i4_3_lut_4_lut (.A(n15018), .B(n15022), .C(\array[251] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_4065[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_8_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_8_i5_3_lut_4_lut (.A(n15018), .B(n15022), .C(\array[251] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_4065[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_8_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_8_i6_3_lut_4_lut (.A(n15018), .B(n15022), .C(\array[251] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_4065[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_8_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_8_i7_3_lut_4_lut (.A(n15018), .B(n15022), .C(\array[251] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_4065[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_8_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_8_i8_3_lut_4_lut (.A(n15018), .B(n15022), .C(\array[251] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_4065[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_8_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_7_i1_3_lut_4_lut (.A(n15019), .B(n15022), .C(\array[252] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_4073[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_7_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_7_i2_3_lut_4_lut (.A(n15019), .B(n15022), .C(\array[252] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_4073[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_7_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_7_i3_3_lut_4_lut (.A(n15019), .B(n15022), .C(\array[252] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_4073[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_7_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_7_i4_3_lut_4_lut (.A(n15019), .B(n15022), .C(\array[252] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_4073[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_7_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_7_i5_3_lut_4_lut (.A(n15019), .B(n15022), .C(\array[252] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_4073[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_7_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_7_i6_3_lut_4_lut (.A(n15019), .B(n15022), .C(\array[252] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_4073[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_7_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_7_i7_3_lut_4_lut (.A(n15019), .B(n15022), .C(\array[252] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_4073[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_7_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_7_i8_3_lut_4_lut (.A(n15019), .B(n15022), .C(\array[252] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_4073[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_7_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_6_i1_3_lut_4_lut (.A(n15020), .B(n15022), .C(\array[253] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_4081[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_6_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_6_i2_3_lut_4_lut (.A(n15020), .B(n15022), .C(\array[253] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_4081[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_6_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_6_i3_3_lut_4_lut (.A(n15020), .B(n15022), .C(\array[253] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_4081[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_6_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_6_i4_3_lut_4_lut (.A(n15020), .B(n15022), .C(\array[253] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_4081[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_6_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_6_i5_3_lut_4_lut (.A(n15020), .B(n15022), .C(\array[253] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_4081[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_6_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_6_i6_3_lut_4_lut (.A(n15020), .B(n15022), .C(\array[253] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_4081[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_6_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_6_i7_3_lut_4_lut (.A(n15020), .B(n15022), .C(\array[253] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_4081[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_6_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_6_i8_3_lut_4_lut (.A(n15020), .B(n15022), .C(\array[253] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_4081[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_6_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_5_i1_3_lut_4_lut (.A(n15021), .B(n15022), .C(\array[254] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_4089[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_5_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_5_i2_3_lut_4_lut (.A(n15021), .B(n15022), .C(\array[254] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_4089[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_5_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_5_i3_3_lut_4_lut (.A(n15021), .B(n15022), .C(\array[254] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_4089[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_5_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_5_i4_3_lut_4_lut (.A(n15021), .B(n15022), .C(\array[254] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_4089[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_5_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_5_i5_3_lut_4_lut (.A(n15021), .B(n15022), .C(\array[254] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_4089[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_5_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_5_i6_3_lut_4_lut (.A(n15021), .B(n15022), .C(\array[254] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_4089[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_5_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_5_i7_3_lut_4_lut (.A(n15021), .B(n15022), .C(\array[254] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_4089[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_5_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_5_i8_3_lut_4_lut (.A(n15021), .B(n15022), .C(\array[254] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_4089[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_5_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_221_i1_3_lut_4_lut (.A(n15013), .B(n14994), .C(\array[38] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_2361[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_221_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_221_i2_3_lut_4_lut (.A(n15013), .B(n14994), .C(\array[38] [1]), 
         .D(d_in_c_1), .Z(array_0__7__N_2361[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_221_i2_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX r_addr_i0_i2 (.D(addr_c_2), .SP(clk_c_enable_2057), .CK(clk_c), 
            .Q(r_addr[2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam r_addr_i0_i2.GSR = "ENABLED";
    FD1P3AX r_addr_i0_i3 (.D(addr_c_3), .SP(clk_c_enable_2057), .CK(clk_c), 
            .Q(r_addr[3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam r_addr_i0_i3.GSR = "ENABLED";
    FD1P3AX r_addr_i0_i4 (.D(addr_c_4), .SP(clk_c_enable_2057), .CK(clk_c), 
            .Q(r_addr[4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam r_addr_i0_i4.GSR = "ENABLED";
    FD1P3AX r_addr_i0_i5 (.D(addr_c_5), .SP(clk_c_enable_2057), .CK(clk_c), 
            .Q(r_addr[5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam r_addr_i0_i5.GSR = "ENABLED";
    FD1P3AX r_addr_i0_i6 (.D(addr_c_6), .SP(clk_c_enable_2057), .CK(clk_c), 
            .Q(r_addr[6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam r_addr_i0_i6.GSR = "ENABLED";
    FD1P3AX r_addr_i0_i7 (.D(addr_c_7), .SP(clk_c_enable_2057), .CK(clk_c), 
            .Q(r_addr[7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam r_addr_i0_i7.GSR = "ENABLED";
    FD1P3AX array_255___i2 (.D(array_0__7__N_4097[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[255] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2.GSR = "ENABLED";
    L6MUX21 i5896 (.D0(n14436), .D1(n14437), .SD(r_addr[7]), .Z(d_out_c_6));
    L6MUX21 i5386 (.D0(n13926), .D1(n13927), .SD(r_addr[7]), .Z(d_out_c_4));
    L6MUX21 i4621 (.D0(n13161), .D1(n13162), .SD(r_addr[7]), .Z(d_out_c_1));
    L6MUX21 i5641 (.D0(n14181), .D1(n14182), .SD(r_addr[7]), .Z(d_out_c_5));
    L6MUX21 i4876 (.D0(n13416), .D1(n13417), .SD(r_addr[7]), .Z(d_out_c_2));
    L6MUX21 i6406 (.D0(n14946), .D1(n14947), .SD(r_addr[7]), .Z(d_out_c_0));
    L6MUX21 i5131 (.D0(n13671), .D1(n13672), .SD(r_addr[7]), .Z(d_out_c_3));
    L6MUX21 i6151 (.D0(n14691), .D1(n14692), .SD(r_addr[7]), .Z(d_out_c_7));
    L6MUX21 i5894 (.D0(n14432), .D1(n14433), .SD(r_addr[6]), .Z(n14436));
    L6MUX21 i5895 (.D0(n14434), .D1(n14435), .SD(r_addr[6]), .Z(n14437));
    L6MUX21 i5384 (.D0(n13922), .D1(n13923), .SD(r_addr[6]), .Z(n13926));
    L6MUX21 i5385 (.D0(n13924), .D1(n13925), .SD(r_addr[6]), .Z(n13927));
    L6MUX21 i4619 (.D0(n13157), .D1(n13158), .SD(r_addr[6]), .Z(n13161));
    L6MUX21 i4620 (.D0(n13159), .D1(n13160), .SD(r_addr[6]), .Z(n13162));
    L6MUX21 i6404 (.D0(n14942), .D1(n14943), .SD(r_addr[6]), .Z(n14946));
    L6MUX21 i5639 (.D0(n14177), .D1(n14178), .SD(r_addr[6]), .Z(n14181));
    L6MUX21 i5640 (.D0(n14179), .D1(n14180), .SD(r_addr[6]), .Z(n14182));
    L6MUX21 i4874 (.D0(n13412), .D1(n13413), .SD(r_addr[6]), .Z(n13416));
    L6MUX21 i4875 (.D0(n13414), .D1(n13415), .SD(r_addr[6]), .Z(n13417));
    L6MUX21 i6405 (.D0(n14944), .D1(n14945), .SD(r_addr[6]), .Z(n14947));
    L6MUX21 i5129 (.D0(n13667), .D1(n13668), .SD(r_addr[6]), .Z(n13671));
    L6MUX21 i5130 (.D0(n13669), .D1(n13670), .SD(r_addr[6]), .Z(n13672));
    L6MUX21 i6149 (.D0(n14687), .D1(n14688), .SD(r_addr[6]), .Z(n14691));
    L6MUX21 i6150 (.D0(n14689), .D1(n14690), .SD(r_addr[6]), .Z(n14692));
    PFUMX i5891 (.BLUT(n14276), .ALUT(n14307), .C0(r_addr[5]), .Z(n14433));
    PFUMX i5892 (.BLUT(n14338), .ALUT(n14369), .C0(r_addr[5]), .Z(n14434));
    PFUMX i5893 (.BLUT(n14400), .ALUT(n14431), .C0(r_addr[5]), .Z(n14435));
    PFUMX i5381 (.BLUT(n13766), .ALUT(n13797), .C0(r_addr[5]), .Z(n13923));
    PFUMX i5382 (.BLUT(n13828), .ALUT(n13859), .C0(r_addr[5]), .Z(n13924));
    PFUMX i5383 (.BLUT(n13890), .ALUT(n13921), .C0(r_addr[5]), .Z(n13925));
    PFUMX i6401 (.BLUT(n14786), .ALUT(n14817), .C0(r_addr[5]), .Z(n14943));
    PFUMX i6400 (.BLUT(n14724), .ALUT(n14755), .C0(r_addr[5]), .Z(n14942));
    PFUMX i6145 (.BLUT(n14469), .ALUT(n14500), .C0(r_addr[5]), .Z(n14687));
    PFUMX i5890 (.BLUT(n14214), .ALUT(n14245), .C0(r_addr[5]), .Z(n14432));
    PFUMX i5635 (.BLUT(n13959), .ALUT(n13990), .C0(r_addr[5]), .Z(n14177));
    PFUMX i5380 (.BLUT(n13704), .ALUT(n13735), .C0(r_addr[5]), .Z(n13922));
    PFUMX i5125 (.BLUT(n13449), .ALUT(n13480), .C0(r_addr[5]), .Z(n13667));
    PFUMX i4870 (.BLUT(n13194), .ALUT(n13225), .C0(r_addr[5]), .Z(n13412));
    PFUMX i4615 (.BLUT(n12939), .ALUT(n12970), .C0(r_addr[5]), .Z(n13157));
    PFUMX i6402 (.BLUT(n14848), .ALUT(n14879), .C0(r_addr[5]), .Z(n14944));
    PFUMX i4616 (.BLUT(n13001), .ALUT(n13032), .C0(r_addr[5]), .Z(n13158));
    PFUMX i4617 (.BLUT(n13063), .ALUT(n13094), .C0(r_addr[5]), .Z(n13159));
    PFUMX i4618 (.BLUT(n13125), .ALUT(n13156), .C0(r_addr[5]), .Z(n13160));
    PFUMX i6403 (.BLUT(n14910), .ALUT(n14941), .C0(r_addr[5]), .Z(n14945));
    PFUMX i5636 (.BLUT(n14021), .ALUT(n14052), .C0(r_addr[5]), .Z(n14178));
    PFUMX i5637 (.BLUT(n14083), .ALUT(n14114), .C0(r_addr[5]), .Z(n14179));
    PFUMX i5638 (.BLUT(n14145), .ALUT(n14176), .C0(r_addr[5]), .Z(n14180));
    PFUMX i4871 (.BLUT(n13256), .ALUT(n13287), .C0(r_addr[5]), .Z(n13413));
    PFUMX i4872 (.BLUT(n13318), .ALUT(n13349), .C0(r_addr[5]), .Z(n13414));
    PFUMX i4873 (.BLUT(n13380), .ALUT(n13411), .C0(r_addr[5]), .Z(n13415));
    PFUMX i5126 (.BLUT(n13511), .ALUT(n13542), .C0(r_addr[5]), .Z(n13668));
    PFUMX i5127 (.BLUT(n13573), .ALUT(n13604), .C0(r_addr[5]), .Z(n13669));
    PFUMX i5128 (.BLUT(n13635), .ALUT(n13666), .C0(r_addr[5]), .Z(n13670));
    PFUMX i6146 (.BLUT(n14531), .ALUT(n14562), .C0(r_addr[5]), .Z(n14688));
    PFUMX i6147 (.BLUT(n14593), .ALUT(n14624), .C0(r_addr[5]), .Z(n14689));
    PFUMX i6148 (.BLUT(n14655), .ALUT(n14686), .C0(r_addr[5]), .Z(n14690));
    L6MUX21 i5887 (.D0(n14425), .D1(n14426), .SD(r_addr[3]), .Z(n14429));
    L6MUX21 i5888 (.D0(n14427), .D1(n14428), .SD(r_addr[3]), .Z(n14430));
    L6MUX21 i4395 (.D0(n12933), .D1(n12934), .SD(r_addr[3]), .Z(n12937));
    L6MUX21 i4396 (.D0(n12935), .D1(n12936), .SD(r_addr[3]), .Z(n12938));
    L6MUX21 i5377 (.D0(n13915), .D1(n13916), .SD(r_addr[3]), .Z(n13919));
    L6MUX21 i5378 (.D0(n13917), .D1(n13918), .SD(r_addr[3]), .Z(n13920));
    L6MUX21 i4426 (.D0(n12964), .D1(n12965), .SD(r_addr[3]), .Z(n12968));
    L6MUX21 i4427 (.D0(n12966), .D1(n12967), .SD(r_addr[3]), .Z(n12969));
    L6MUX21 i4457 (.D0(n12995), .D1(n12996), .SD(r_addr[3]), .Z(n12999));
    L6MUX21 i4458 (.D0(n12997), .D1(n12998), .SD(r_addr[3]), .Z(n13000));
    L6MUX21 i4488 (.D0(n13026), .D1(n13027), .SD(r_addr[3]), .Z(n13030));
    L6MUX21 i5415 (.D0(n13953), .D1(n13954), .SD(r_addr[3]), .Z(n13957));
    L6MUX21 i4489 (.D0(n13028), .D1(n13029), .SD(r_addr[3]), .Z(n13031));
    L6MUX21 i5416 (.D0(n13955), .D1(n13956), .SD(r_addr[3]), .Z(n13958));
    L6MUX21 i4519 (.D0(n13057), .D1(n13058), .SD(r_addr[3]), .Z(n13061));
    L6MUX21 i4520 (.D0(n13059), .D1(n13060), .SD(r_addr[3]), .Z(n13062));
    L6MUX21 i5925 (.D0(n14463), .D1(n14464), .SD(r_addr[3]), .Z(n14467));
    L6MUX21 i5926 (.D0(n14465), .D1(n14466), .SD(r_addr[3]), .Z(n14468));
    L6MUX21 i5446 (.D0(n13984), .D1(n13985), .SD(r_addr[3]), .Z(n13988));
    L6MUX21 i5447 (.D0(n13986), .D1(n13987), .SD(r_addr[3]), .Z(n13989));
    L6MUX21 i6180 (.D0(n14718), .D1(n14719), .SD(r_addr[3]), .Z(n14722));
    L6MUX21 i5477 (.D0(n14015), .D1(n14016), .SD(r_addr[3]), .Z(n14019));
    L6MUX21 i6181 (.D0(n14720), .D1(n14721), .SD(r_addr[3]), .Z(n14723));
    L6MUX21 i5478 (.D0(n14017), .D1(n14018), .SD(r_addr[3]), .Z(n14020));
    L6MUX21 i4550 (.D0(n13088), .D1(n13089), .SD(r_addr[3]), .Z(n13092));
    L6MUX21 i4551 (.D0(n13090), .D1(n13091), .SD(r_addr[3]), .Z(n13093));
    L6MUX21 i5956 (.D0(n14494), .D1(n14495), .SD(r_addr[3]), .Z(n14498));
    L6MUX21 i5957 (.D0(n14496), .D1(n14497), .SD(r_addr[3]), .Z(n14499));
    L6MUX21 i4581 (.D0(n13119), .D1(n13120), .SD(r_addr[3]), .Z(n13123));
    L6MUX21 i4582 (.D0(n13121), .D1(n13122), .SD(r_addr[3]), .Z(n13124));
    L6MUX21 i5508 (.D0(n14046), .D1(n14047), .SD(r_addr[3]), .Z(n14050));
    L6MUX21 i5509 (.D0(n14048), .D1(n14049), .SD(r_addr[3]), .Z(n14051));
    L6MUX21 i4612 (.D0(n13150), .D1(n13151), .SD(r_addr[3]), .Z(n13154));
    L6MUX21 i4613 (.D0(n13152), .D1(n13153), .SD(r_addr[3]), .Z(n13155));
    L6MUX21 i6304 (.D0(n14842), .D1(n14843), .SD(r_addr[3]), .Z(n14846));
    L6MUX21 i6305 (.D0(n14844), .D1(n14845), .SD(r_addr[3]), .Z(n14847));
    L6MUX21 i4650 (.D0(n13188), .D1(n13189), .SD(r_addr[3]), .Z(n13192));
    L6MUX21 i4651 (.D0(n13190), .D1(n13191), .SD(r_addr[3]), .Z(n13193));
    L6MUX21 i5539 (.D0(n14077), .D1(n14078), .SD(r_addr[3]), .Z(n14081));
    L6MUX21 i5540 (.D0(n14079), .D1(n14080), .SD(r_addr[3]), .Z(n14082));
    L6MUX21 i4681 (.D0(n13219), .D1(n13220), .SD(r_addr[3]), .Z(n13223));
    L6MUX21 i4682 (.D0(n13221), .D1(n13222), .SD(r_addr[3]), .Z(n13224));
    L6MUX21 i5987 (.D0(n14525), .D1(n14526), .SD(r_addr[3]), .Z(n14529));
    L6MUX21 i5988 (.D0(n14527), .D1(n14528), .SD(r_addr[3]), .Z(n14530));
    L6MUX21 i4712 (.D0(n13250), .D1(n13251), .SD(r_addr[3]), .Z(n13254));
    L6MUX21 i4713 (.D0(n13252), .D1(n13253), .SD(r_addr[3]), .Z(n13255));
    L6MUX21 i5570 (.D0(n14108), .D1(n14109), .SD(r_addr[3]), .Z(n14112));
    L6MUX21 i5571 (.D0(n14110), .D1(n14111), .SD(r_addr[3]), .Z(n14113));
    L6MUX21 i4743 (.D0(n13281), .D1(n13282), .SD(r_addr[3]), .Z(n13285));
    L6MUX21 i4744 (.D0(n13283), .D1(n13284), .SD(r_addr[3]), .Z(n13286));
    L6MUX21 i4774 (.D0(n13312), .D1(n13313), .SD(r_addr[3]), .Z(n13316));
    L6MUX21 i4775 (.D0(n13314), .D1(n13315), .SD(r_addr[3]), .Z(n13317));
    L6MUX21 i6211 (.D0(n14749), .D1(n14750), .SD(r_addr[3]), .Z(n14753));
    L6MUX21 i5601 (.D0(n14139), .D1(n14140), .SD(r_addr[3]), .Z(n14143));
    L6MUX21 i6212 (.D0(n14751), .D1(n14752), .SD(r_addr[3]), .Z(n14754));
    L6MUX21 i5602 (.D0(n14141), .D1(n14142), .SD(r_addr[3]), .Z(n14144));
    L6MUX21 i4805 (.D0(n13343), .D1(n13344), .SD(r_addr[3]), .Z(n13347));
    L6MUX21 i4806 (.D0(n13345), .D1(n13346), .SD(r_addr[3]), .Z(n13348));
    L6MUX21 i6018 (.D0(n14556), .D1(n14557), .SD(r_addr[3]), .Z(n14560));
    L6MUX21 i6366 (.D0(n14904), .D1(n14905), .SD(r_addr[3]), .Z(n14908));
    L6MUX21 i6019 (.D0(n14558), .D1(n14559), .SD(r_addr[3]), .Z(n14561));
    L6MUX21 i4836 (.D0(n13374), .D1(n13375), .SD(r_addr[3]), .Z(n13378));
    L6MUX21 i4837 (.D0(n13376), .D1(n13377), .SD(r_addr[3]), .Z(n13379));
    L6MUX21 i5632 (.D0(n14170), .D1(n14171), .SD(r_addr[3]), .Z(n14174));
    L6MUX21 i5633 (.D0(n14172), .D1(n14173), .SD(r_addr[3]), .Z(n14175));
    L6MUX21 i6367 (.D0(n14906), .D1(n14907), .SD(r_addr[3]), .Z(n14909));
    L6MUX21 i4867 (.D0(n13405), .D1(n13406), .SD(r_addr[3]), .Z(n13409));
    L6MUX21 i4868 (.D0(n13407), .D1(n13408), .SD(r_addr[3]), .Z(n13410));
    L6MUX21 i4905 (.D0(n13443), .D1(n13444), .SD(r_addr[3]), .Z(n13447));
    L6MUX21 i4906 (.D0(n13445), .D1(n13446), .SD(r_addr[3]), .Z(n13448));
    L6MUX21 i5670 (.D0(n14208), .D1(n14209), .SD(r_addr[3]), .Z(n14212));
    L6MUX21 i5671 (.D0(n14210), .D1(n14211), .SD(r_addr[3]), .Z(n14213));
    L6MUX21 i4936 (.D0(n13474), .D1(n13475), .SD(r_addr[3]), .Z(n13478));
    L6MUX21 i4937 (.D0(n13476), .D1(n13477), .SD(r_addr[3]), .Z(n13479));
    L6MUX21 i6049 (.D0(n14587), .D1(n14588), .SD(r_addr[3]), .Z(n14591));
    L6MUX21 i6050 (.D0(n14589), .D1(n14590), .SD(r_addr[3]), .Z(n14592));
    L6MUX21 i4967 (.D0(n13505), .D1(n13506), .SD(r_addr[3]), .Z(n13509));
    L6MUX21 i4968 (.D0(n13507), .D1(n13508), .SD(r_addr[3]), .Z(n13510));
    L6MUX21 i5701 (.D0(n14239), .D1(n14240), .SD(r_addr[3]), .Z(n14243));
    L6MUX21 i5702 (.D0(n14241), .D1(n14242), .SD(r_addr[3]), .Z(n14244));
    L6MUX21 i4998 (.D0(n13536), .D1(n13537), .SD(r_addr[3]), .Z(n13540));
    L6MUX21 i4999 (.D0(n13538), .D1(n13539), .SD(r_addr[3]), .Z(n13541));
    L6MUX21 i6242 (.D0(n14780), .D1(n14781), .SD(r_addr[3]), .Z(n14784));
    L6MUX21 i5029 (.D0(n13567), .D1(n13568), .SD(r_addr[3]), .Z(n13571));
    L6MUX21 i5030 (.D0(n13569), .D1(n13570), .SD(r_addr[3]), .Z(n13572));
    L6MUX21 i6243 (.D0(n14782), .D1(n14783), .SD(r_addr[3]), .Z(n14785));
    L6MUX21 i5732 (.D0(n14270), .D1(n14271), .SD(r_addr[3]), .Z(n14274));
    L6MUX21 i5733 (.D0(n14272), .D1(n14273), .SD(r_addr[3]), .Z(n14275));
    L6MUX21 i5060 (.D0(n13598), .D1(n13599), .SD(r_addr[3]), .Z(n13602));
    L6MUX21 i5061 (.D0(n13600), .D1(n13601), .SD(r_addr[3]), .Z(n13603));
    L6MUX21 i6080 (.D0(n14618), .D1(n14619), .SD(r_addr[3]), .Z(n14622));
    L6MUX21 i6081 (.D0(n14620), .D1(n14621), .SD(r_addr[3]), .Z(n14623));
    L6MUX21 i5091 (.D0(n13629), .D1(n13630), .SD(r_addr[3]), .Z(n13633));
    L6MUX21 i5092 (.D0(n13631), .D1(n13632), .SD(r_addr[3]), .Z(n13634));
    L6MUX21 i5763 (.D0(n14301), .D1(n14302), .SD(r_addr[3]), .Z(n14305));
    L6MUX21 i5764 (.D0(n14303), .D1(n14304), .SD(r_addr[3]), .Z(n14306));
    L6MUX21 i6335 (.D0(n14873), .D1(n14874), .SD(r_addr[3]), .Z(n14877));
    L6MUX21 i5122 (.D0(n13660), .D1(n13661), .SD(r_addr[3]), .Z(n13664));
    L6MUX21 i5123 (.D0(n13662), .D1(n13663), .SD(r_addr[3]), .Z(n13665));
    L6MUX21 i6336 (.D0(n14875), .D1(n14876), .SD(r_addr[3]), .Z(n14878));
    L6MUX21 i5160 (.D0(n13698), .D1(n13699), .SD(r_addr[3]), .Z(n13702));
    L6MUX21 i5161 (.D0(n13700), .D1(n13701), .SD(r_addr[3]), .Z(n13703));
    L6MUX21 i5794 (.D0(n14332), .D1(n14333), .SD(r_addr[3]), .Z(n14336));
    L6MUX21 i5795 (.D0(n14334), .D1(n14335), .SD(r_addr[3]), .Z(n14337));
    L6MUX21 i6111 (.D0(n14649), .D1(n14650), .SD(r_addr[3]), .Z(n14653));
    L6MUX21 i5191 (.D0(n13729), .D1(n13730), .SD(r_addr[3]), .Z(n13733));
    L6MUX21 i5192 (.D0(n13731), .D1(n13732), .SD(r_addr[3]), .Z(n13734));
    L6MUX21 i6112 (.D0(n14651), .D1(n14652), .SD(r_addr[3]), .Z(n14654));
    L6MUX21 i6397 (.D0(n14935), .D1(n14936), .SD(r_addr[3]), .Z(n14939));
    L6MUX21 i5222 (.D0(n13760), .D1(n13761), .SD(r_addr[3]), .Z(n13764));
    L6MUX21 i5223 (.D0(n13762), .D1(n13763), .SD(r_addr[3]), .Z(n13765));
    L6MUX21 i5825 (.D0(n14363), .D1(n14364), .SD(r_addr[3]), .Z(n14367));
    L6MUX21 i5826 (.D0(n14365), .D1(n14366), .SD(r_addr[3]), .Z(n14368));
    L6MUX21 i5253 (.D0(n13791), .D1(n13792), .SD(r_addr[3]), .Z(n13795));
    L6MUX21 i5254 (.D0(n13793), .D1(n13794), .SD(r_addr[3]), .Z(n13796));
    L6MUX21 i6273 (.D0(n14811), .D1(n14812), .SD(r_addr[3]), .Z(n14815));
    L6MUX21 i6274 (.D0(n14813), .D1(n14814), .SD(r_addr[3]), .Z(n14816));
    L6MUX21 i5284 (.D0(n13822), .D1(n13823), .SD(r_addr[3]), .Z(n13826));
    L6MUX21 i6398 (.D0(n14937), .D1(n14938), .SD(r_addr[3]), .Z(n14940));
    L6MUX21 i5285 (.D0(n13824), .D1(n13825), .SD(r_addr[3]), .Z(n13827));
    L6MUX21 i5856 (.D0(n14394), .D1(n14395), .SD(r_addr[3]), .Z(n14398));
    L6MUX21 i5857 (.D0(n14396), .D1(n14397), .SD(r_addr[3]), .Z(n14399));
    L6MUX21 i6142 (.D0(n14680), .D1(n14681), .SD(r_addr[3]), .Z(n14684));
    L6MUX21 i5315 (.D0(n13853), .D1(n13854), .SD(r_addr[3]), .Z(n13857));
    L6MUX21 i5316 (.D0(n13855), .D1(n13856), .SD(r_addr[3]), .Z(n13858));
    L6MUX21 i6143 (.D0(n14682), .D1(n14683), .SD(r_addr[3]), .Z(n14685));
    L6MUX21 i5346 (.D0(n13884), .D1(n13885), .SD(r_addr[3]), .Z(n13888));
    L6MUX21 i5347 (.D0(n13886), .D1(n13887), .SD(r_addr[3]), .Z(n13889));
    L6MUX21 i4391 (.D0(n12925), .D1(n12926), .SD(r_addr[2]), .Z(n12933));
    L6MUX21 i4392 (.D0(n12927), .D1(n12928), .SD(r_addr[2]), .Z(n12934));
    L6MUX21 i4393 (.D0(n12929), .D1(n12930), .SD(r_addr[2]), .Z(n12935));
    L6MUX21 i4394 (.D0(n12931), .D1(n12932), .SD(r_addr[2]), .Z(n12936));
    L6MUX21 i5373 (.D0(n13907), .D1(n13908), .SD(r_addr[2]), .Z(n13915));
    L6MUX21 i5374 (.D0(n13909), .D1(n13910), .SD(r_addr[2]), .Z(n13916));
    L6MUX21 i5375 (.D0(n13911), .D1(n13912), .SD(r_addr[2]), .Z(n13917));
    L6MUX21 i5376 (.D0(n13913), .D1(n13914), .SD(r_addr[2]), .Z(n13918));
    L6MUX21 i4422 (.D0(n12956), .D1(n12957), .SD(r_addr[2]), .Z(n12964));
    L6MUX21 i4423 (.D0(n12958), .D1(n12959), .SD(r_addr[2]), .Z(n12965));
    L6MUX21 i4424 (.D0(n12960), .D1(n12961), .SD(r_addr[2]), .Z(n12966));
    L6MUX21 i4425 (.D0(n12962), .D1(n12963), .SD(r_addr[2]), .Z(n12967));
    L6MUX21 i4453 (.D0(n12987), .D1(n12988), .SD(r_addr[2]), .Z(n12995));
    L6MUX21 i4454 (.D0(n12989), .D1(n12990), .SD(r_addr[2]), .Z(n12996));
    L6MUX21 i4455 (.D0(n12991), .D1(n12992), .SD(r_addr[2]), .Z(n12997));
    L6MUX21 i4456 (.D0(n12993), .D1(n12994), .SD(r_addr[2]), .Z(n12998));
    L6MUX21 i5411 (.D0(n13945), .D1(n13946), .SD(r_addr[2]), .Z(n13953));
    L6MUX21 i5412 (.D0(n13947), .D1(n13948), .SD(r_addr[2]), .Z(n13954));
    L6MUX21 i4484 (.D0(n13018), .D1(n13019), .SD(r_addr[2]), .Z(n13026));
    L6MUX21 i5413 (.D0(n13949), .D1(n13950), .SD(r_addr[2]), .Z(n13955));
    L6MUX21 i4485 (.D0(n13020), .D1(n13021), .SD(r_addr[2]), .Z(n13027));
    L6MUX21 i4486 (.D0(n13022), .D1(n13023), .SD(r_addr[2]), .Z(n13028));
    L6MUX21 i5414 (.D0(n13951), .D1(n13952), .SD(r_addr[2]), .Z(n13956));
    L6MUX21 i4487 (.D0(n13024), .D1(n13025), .SD(r_addr[2]), .Z(n13029));
    L6MUX21 i5921 (.D0(n14455), .D1(n14456), .SD(r_addr[2]), .Z(n14463));
    L6MUX21 i5922 (.D0(n14457), .D1(n14458), .SD(r_addr[2]), .Z(n14464));
    L6MUX21 i4515 (.D0(n13049), .D1(n13050), .SD(r_addr[2]), .Z(n13057));
    L6MUX21 i4516 (.D0(n13051), .D1(n13052), .SD(r_addr[2]), .Z(n13058));
    L6MUX21 i4517 (.D0(n13053), .D1(n13054), .SD(r_addr[2]), .Z(n13059));
    L6MUX21 i4518 (.D0(n13055), .D1(n13056), .SD(r_addr[2]), .Z(n13060));
    L6MUX21 i5923 (.D0(n14459), .D1(n14460), .SD(r_addr[2]), .Z(n14465));
    L6MUX21 i5924 (.D0(n14461), .D1(n14462), .SD(r_addr[2]), .Z(n14466));
    L6MUX21 i5442 (.D0(n13976), .D1(n13977), .SD(r_addr[2]), .Z(n13984));
    L6MUX21 i5443 (.D0(n13978), .D1(n13979), .SD(r_addr[2]), .Z(n13985));
    L6MUX21 i5444 (.D0(n13980), .D1(n13981), .SD(r_addr[2]), .Z(n13986));
    L6MUX21 i5445 (.D0(n13982), .D1(n13983), .SD(r_addr[2]), .Z(n13987));
    L6MUX21 i6176 (.D0(n14710), .D1(n14711), .SD(r_addr[2]), .Z(n14718));
    L6MUX21 i6177 (.D0(n14712), .D1(n14713), .SD(r_addr[2]), .Z(n14719));
    L6MUX21 i6178 (.D0(n14714), .D1(n14715), .SD(r_addr[2]), .Z(n14720));
    L6MUX21 i6179 (.D0(n14716), .D1(n14717), .SD(r_addr[2]), .Z(n14721));
    L6MUX21 i5473 (.D0(n14007), .D1(n14008), .SD(r_addr[2]), .Z(n14015));
    L6MUX21 i5474 (.D0(n14009), .D1(n14010), .SD(r_addr[2]), .Z(n14016));
    L6MUX21 i5475 (.D0(n14011), .D1(n14012), .SD(r_addr[2]), .Z(n14017));
    L6MUX21 i5476 (.D0(n14013), .D1(n14014), .SD(r_addr[2]), .Z(n14018));
    L6MUX21 i4546 (.D0(n13080), .D1(n13081), .SD(r_addr[2]), .Z(n13088));
    L6MUX21 i4547 (.D0(n13082), .D1(n13083), .SD(r_addr[2]), .Z(n13089));
    L6MUX21 i4548 (.D0(n13084), .D1(n13085), .SD(r_addr[2]), .Z(n13090));
    L6MUX21 i4549 (.D0(n13086), .D1(n13087), .SD(r_addr[2]), .Z(n13091));
    L6MUX21 i5952 (.D0(n14486), .D1(n14487), .SD(r_addr[2]), .Z(n14494));
    L6MUX21 i6300 (.D0(n14834), .D1(n14835), .SD(r_addr[2]), .Z(n14842));
    L6MUX21 i5953 (.D0(n14488), .D1(n14489), .SD(r_addr[2]), .Z(n14495));
    L6MUX21 i5954 (.D0(n14490), .D1(n14491), .SD(r_addr[2]), .Z(n14496));
    L6MUX21 i5955 (.D0(n14492), .D1(n14493), .SD(r_addr[2]), .Z(n14497));
    L6MUX21 i4577 (.D0(n13111), .D1(n13112), .SD(r_addr[2]), .Z(n13119));
    L6MUX21 i4578 (.D0(n13113), .D1(n13114), .SD(r_addr[2]), .Z(n13120));
    L6MUX21 i4579 (.D0(n13115), .D1(n13116), .SD(r_addr[2]), .Z(n13121));
    L6MUX21 i6301 (.D0(n14836), .D1(n14837), .SD(r_addr[2]), .Z(n14843));
    L6MUX21 i4580 (.D0(n13117), .D1(n13118), .SD(r_addr[2]), .Z(n13122));
    L6MUX21 i5504 (.D0(n14038), .D1(n14039), .SD(r_addr[2]), .Z(n14046));
    L6MUX21 i5505 (.D0(n14040), .D1(n14041), .SD(r_addr[2]), .Z(n14047));
    L6MUX21 i5506 (.D0(n14042), .D1(n14043), .SD(r_addr[2]), .Z(n14048));
    L6MUX21 i6302 (.D0(n14838), .D1(n14839), .SD(r_addr[2]), .Z(n14844));
    L6MUX21 i5507 (.D0(n14044), .D1(n14045), .SD(r_addr[2]), .Z(n14049));
    L6MUX21 i4608 (.D0(n13142), .D1(n13143), .SD(r_addr[2]), .Z(n13150));
    L6MUX21 i4609 (.D0(n13144), .D1(n13145), .SD(r_addr[2]), .Z(n13151));
    L6MUX21 i4610 (.D0(n13146), .D1(n13147), .SD(r_addr[2]), .Z(n13152));
    L6MUX21 i4611 (.D0(n13148), .D1(n13149), .SD(r_addr[2]), .Z(n13153));
    L6MUX21 i6303 (.D0(n14840), .D1(n14841), .SD(r_addr[2]), .Z(n14845));
    L6MUX21 i4646 (.D0(n13180), .D1(n13181), .SD(r_addr[2]), .Z(n13188));
    L6MUX21 i4647 (.D0(n13182), .D1(n13183), .SD(r_addr[2]), .Z(n13189));
    L6MUX21 i4648 (.D0(n13184), .D1(n13185), .SD(r_addr[2]), .Z(n13190));
    L6MUX21 i4649 (.D0(n13186), .D1(n13187), .SD(r_addr[2]), .Z(n13191));
    L6MUX21 i5535 (.D0(n14069), .D1(n14070), .SD(r_addr[2]), .Z(n14077));
    L6MUX21 i5536 (.D0(n14071), .D1(n14072), .SD(r_addr[2]), .Z(n14078));
    L6MUX21 i5537 (.D0(n14073), .D1(n14074), .SD(r_addr[2]), .Z(n14079));
    L6MUX21 i5538 (.D0(n14075), .D1(n14076), .SD(r_addr[2]), .Z(n14080));
    L6MUX21 i4677 (.D0(n13211), .D1(n13212), .SD(r_addr[2]), .Z(n13219));
    L6MUX21 i4678 (.D0(n13213), .D1(n13214), .SD(r_addr[2]), .Z(n13220));
    L6MUX21 i4679 (.D0(n13215), .D1(n13216), .SD(r_addr[2]), .Z(n13221));
    L6MUX21 i4680 (.D0(n13217), .D1(n13218), .SD(r_addr[2]), .Z(n13222));
    L6MUX21 i5983 (.D0(n14517), .D1(n14518), .SD(r_addr[2]), .Z(n14525));
    L6MUX21 i5984 (.D0(n14519), .D1(n14520), .SD(r_addr[2]), .Z(n14526));
    L6MUX21 i5985 (.D0(n14521), .D1(n14522), .SD(r_addr[2]), .Z(n14527));
    L6MUX21 i6362 (.D0(n14896), .D1(n14897), .SD(r_addr[2]), .Z(n14904));
    L6MUX21 i5986 (.D0(n14523), .D1(n14524), .SD(r_addr[2]), .Z(n14528));
    L6MUX21 i4708 (.D0(n13242), .D1(n13243), .SD(r_addr[2]), .Z(n13250));
    L6MUX21 i4709 (.D0(n13244), .D1(n13245), .SD(r_addr[2]), .Z(n13251));
    L6MUX21 i4710 (.D0(n13246), .D1(n13247), .SD(r_addr[2]), .Z(n13252));
    L6MUX21 i4711 (.D0(n13248), .D1(n13249), .SD(r_addr[2]), .Z(n13253));
    L6MUX21 i5566 (.D0(n14100), .D1(n14101), .SD(r_addr[2]), .Z(n14108));
    L6MUX21 i5567 (.D0(n14102), .D1(n14103), .SD(r_addr[2]), .Z(n14109));
    L6MUX21 i5568 (.D0(n14104), .D1(n14105), .SD(r_addr[2]), .Z(n14110));
    L6MUX21 i5569 (.D0(n14106), .D1(n14107), .SD(r_addr[2]), .Z(n14111));
    L6MUX21 i6363 (.D0(n14898), .D1(n14899), .SD(r_addr[2]), .Z(n14905));
    L6MUX21 i4739 (.D0(n13273), .D1(n13274), .SD(r_addr[2]), .Z(n13281));
    L6MUX21 i4740 (.D0(n13275), .D1(n13276), .SD(r_addr[2]), .Z(n13282));
    L6MUX21 i4741 (.D0(n13277), .D1(n13278), .SD(r_addr[2]), .Z(n13283));
    L6MUX21 i4742 (.D0(n13279), .D1(n13280), .SD(r_addr[2]), .Z(n13284));
    L6MUX21 i6207 (.D0(n14741), .D1(n14742), .SD(r_addr[2]), .Z(n14749));
    L6MUX21 i6208 (.D0(n14743), .D1(n14744), .SD(r_addr[2]), .Z(n14750));
    L6MUX21 i6364 (.D0(n14900), .D1(n14901), .SD(r_addr[2]), .Z(n14906));
    L6MUX21 i6209 (.D0(n14745), .D1(n14746), .SD(r_addr[2]), .Z(n14751));
    L6MUX21 i6210 (.D0(n14747), .D1(n14748), .SD(r_addr[2]), .Z(n14752));
    L6MUX21 i4770 (.D0(n13304), .D1(n13305), .SD(r_addr[2]), .Z(n13312));
    L6MUX21 i4771 (.D0(n13306), .D1(n13307), .SD(r_addr[2]), .Z(n13313));
    L6MUX21 i4772 (.D0(n13308), .D1(n13309), .SD(r_addr[2]), .Z(n13314));
    L6MUX21 i4773 (.D0(n13310), .D1(n13311), .SD(r_addr[2]), .Z(n13315));
    L6MUX21 i5597 (.D0(n14131), .D1(n14132), .SD(r_addr[2]), .Z(n14139));
    L6MUX21 i5598 (.D0(n14133), .D1(n14134), .SD(r_addr[2]), .Z(n14140));
    L6MUX21 i5599 (.D0(n14135), .D1(n14136), .SD(r_addr[2]), .Z(n14141));
    L6MUX21 i5600 (.D0(n14137), .D1(n14138), .SD(r_addr[2]), .Z(n14142));
    L6MUX21 i6365 (.D0(n14902), .D1(n14903), .SD(r_addr[2]), .Z(n14907));
    L6MUX21 i4801 (.D0(n13335), .D1(n13336), .SD(r_addr[2]), .Z(n13343));
    L6MUX21 i4802 (.D0(n13337), .D1(n13338), .SD(r_addr[2]), .Z(n13344));
    L6MUX21 i4803 (.D0(n13339), .D1(n13340), .SD(r_addr[2]), .Z(n13345));
    L6MUX21 i4804 (.D0(n13341), .D1(n13342), .SD(r_addr[2]), .Z(n13346));
    L6MUX21 i6014 (.D0(n14548), .D1(n14549), .SD(r_addr[2]), .Z(n14556));
    L6MUX21 i6015 (.D0(n14550), .D1(n14551), .SD(r_addr[2]), .Z(n14557));
    L6MUX21 i6016 (.D0(n14552), .D1(n14553), .SD(r_addr[2]), .Z(n14558));
    L6MUX21 i6017 (.D0(n14554), .D1(n14555), .SD(r_addr[2]), .Z(n14559));
    L6MUX21 i4832 (.D0(n13366), .D1(n13367), .SD(r_addr[2]), .Z(n13374));
    L6MUX21 i4833 (.D0(n13368), .D1(n13369), .SD(r_addr[2]), .Z(n13375));
    L6MUX21 i4834 (.D0(n13370), .D1(n13371), .SD(r_addr[2]), .Z(n13376));
    L6MUX21 i4835 (.D0(n13372), .D1(n13373), .SD(r_addr[2]), .Z(n13377));
    L6MUX21 i5628 (.D0(n14162), .D1(n14163), .SD(r_addr[2]), .Z(n14170));
    L6MUX21 i5629 (.D0(n14164), .D1(n14165), .SD(r_addr[2]), .Z(n14171));
    L6MUX21 i5630 (.D0(n14166), .D1(n14167), .SD(r_addr[2]), .Z(n14172));
    L6MUX21 i5631 (.D0(n14168), .D1(n14169), .SD(r_addr[2]), .Z(n14173));
    L6MUX21 i4863 (.D0(n13397), .D1(n13398), .SD(r_addr[2]), .Z(n13405));
    L6MUX21 i4864 (.D0(n13399), .D1(n13400), .SD(r_addr[2]), .Z(n13406));
    L6MUX21 i4865 (.D0(n13401), .D1(n13402), .SD(r_addr[2]), .Z(n13407));
    L6MUX21 i4866 (.D0(n13403), .D1(n13404), .SD(r_addr[2]), .Z(n13408));
    L6MUX21 i4901 (.D0(n13435), .D1(n13436), .SD(r_addr[2]), .Z(n13443));
    L6MUX21 i4902 (.D0(n13437), .D1(n13438), .SD(r_addr[2]), .Z(n13444));
    L6MUX21 i4903 (.D0(n13439), .D1(n13440), .SD(r_addr[2]), .Z(n13445));
    L6MUX21 i4904 (.D0(n13441), .D1(n13442), .SD(r_addr[2]), .Z(n13446));
    L6MUX21 i5666 (.D0(n14200), .D1(n14201), .SD(r_addr[2]), .Z(n14208));
    L6MUX21 i5667 (.D0(n14202), .D1(n14203), .SD(r_addr[2]), .Z(n14209));
    L6MUX21 i5668 (.D0(n14204), .D1(n14205), .SD(r_addr[2]), .Z(n14210));
    L6MUX21 i5669 (.D0(n14206), .D1(n14207), .SD(r_addr[2]), .Z(n14211));
    L6MUX21 i6045 (.D0(n14579), .D1(n14580), .SD(r_addr[2]), .Z(n14587));
    L6MUX21 i4932 (.D0(n13466), .D1(n13467), .SD(r_addr[2]), .Z(n13474));
    L6MUX21 i6046 (.D0(n14581), .D1(n14582), .SD(r_addr[2]), .Z(n14588));
    L6MUX21 i4933 (.D0(n13468), .D1(n13469), .SD(r_addr[2]), .Z(n13475));
    L6MUX21 i4934 (.D0(n13470), .D1(n13471), .SD(r_addr[2]), .Z(n13476));
    L6MUX21 i4935 (.D0(n13472), .D1(n13473), .SD(r_addr[2]), .Z(n13477));
    L6MUX21 i6047 (.D0(n14583), .D1(n14584), .SD(r_addr[2]), .Z(n14589));
    L6MUX21 i6048 (.D0(n14585), .D1(n14586), .SD(r_addr[2]), .Z(n14590));
    L6MUX21 i6393 (.D0(n14927), .D1(n14928), .SD(r_addr[2]), .Z(n14935));
    L6MUX21 i4963 (.D0(n13497), .D1(n13498), .SD(r_addr[2]), .Z(n13505));
    L6MUX21 i4964 (.D0(n13499), .D1(n13500), .SD(r_addr[2]), .Z(n13506));
    L6MUX21 i4965 (.D0(n13501), .D1(n13502), .SD(r_addr[2]), .Z(n13507));
    L6MUX21 i4966 (.D0(n13503), .D1(n13504), .SD(r_addr[2]), .Z(n13508));
    L6MUX21 i5697 (.D0(n14231), .D1(n14232), .SD(r_addr[2]), .Z(n14239));
    L6MUX21 i5698 (.D0(n14233), .D1(n14234), .SD(r_addr[2]), .Z(n14240));
    L6MUX21 i5699 (.D0(n14235), .D1(n14236), .SD(r_addr[2]), .Z(n14241));
    L6MUX21 i5700 (.D0(n14237), .D1(n14238), .SD(r_addr[2]), .Z(n14242));
    L6MUX21 i6238 (.D0(n14772), .D1(n14773), .SD(r_addr[2]), .Z(n14780));
    L6MUX21 i4994 (.D0(n13528), .D1(n13529), .SD(r_addr[2]), .Z(n13536));
    L6MUX21 i4995 (.D0(n13530), .D1(n13531), .SD(r_addr[2]), .Z(n13537));
    L6MUX21 i4996 (.D0(n13532), .D1(n13533), .SD(r_addr[2]), .Z(n13538));
    L6MUX21 i4997 (.D0(n13534), .D1(n13535), .SD(r_addr[2]), .Z(n13539));
    L6MUX21 i6239 (.D0(n14774), .D1(n14775), .SD(r_addr[2]), .Z(n14781));
    L6MUX21 i6240 (.D0(n14776), .D1(n14777), .SD(r_addr[2]), .Z(n14782));
    L6MUX21 i6241 (.D0(n14778), .D1(n14779), .SD(r_addr[2]), .Z(n14783));
    L6MUX21 i6394 (.D0(n14929), .D1(n14930), .SD(r_addr[2]), .Z(n14936));
    L6MUX21 i5025 (.D0(n13559), .D1(n13560), .SD(r_addr[2]), .Z(n13567));
    L6MUX21 i5026 (.D0(n13561), .D1(n13562), .SD(r_addr[2]), .Z(n13568));
    L6MUX21 i5027 (.D0(n13563), .D1(n13564), .SD(r_addr[2]), .Z(n13569));
    L6MUX21 i5028 (.D0(n13565), .D1(n13566), .SD(r_addr[2]), .Z(n13570));
    L6MUX21 i5728 (.D0(n14262), .D1(n14263), .SD(r_addr[2]), .Z(n14270));
    L6MUX21 i5729 (.D0(n14264), .D1(n14265), .SD(r_addr[2]), .Z(n14271));
    L6MUX21 i5730 (.D0(n14266), .D1(n14267), .SD(r_addr[2]), .Z(n14272));
    L6MUX21 i5731 (.D0(n14268), .D1(n14269), .SD(r_addr[2]), .Z(n14273));
    L6MUX21 i6076 (.D0(n14610), .D1(n14611), .SD(r_addr[2]), .Z(n14618));
    L6MUX21 i6331 (.D0(n14865), .D1(n14866), .SD(r_addr[2]), .Z(n14873));
    L6MUX21 i6077 (.D0(n14612), .D1(n14613), .SD(r_addr[2]), .Z(n14619));
    L6MUX21 i5056 (.D0(n13590), .D1(n13591), .SD(r_addr[2]), .Z(n13598));
    L6MUX21 i5057 (.D0(n13592), .D1(n13593), .SD(r_addr[2]), .Z(n13599));
    L6MUX21 i5058 (.D0(n13594), .D1(n13595), .SD(r_addr[2]), .Z(n13600));
    L6MUX21 i5059 (.D0(n13596), .D1(n13597), .SD(r_addr[2]), .Z(n13601));
    L6MUX21 i6078 (.D0(n14614), .D1(n14615), .SD(r_addr[2]), .Z(n14620));
    L6MUX21 i6079 (.D0(n14616), .D1(n14617), .SD(r_addr[2]), .Z(n14621));
    L6MUX21 i6332 (.D0(n14867), .D1(n14868), .SD(r_addr[2]), .Z(n14874));
    L6MUX21 i5087 (.D0(n13621), .D1(n13622), .SD(r_addr[2]), .Z(n13629));
    L6MUX21 i6395 (.D0(n14931), .D1(n14932), .SD(r_addr[2]), .Z(n14937));
    L6MUX21 i6333 (.D0(n14869), .D1(n14870), .SD(r_addr[2]), .Z(n14875));
    L6MUX21 i5088 (.D0(n13623), .D1(n13624), .SD(r_addr[2]), .Z(n13630));
    L6MUX21 i5089 (.D0(n13625), .D1(n13626), .SD(r_addr[2]), .Z(n13631));
    L6MUX21 i5090 (.D0(n13627), .D1(n13628), .SD(r_addr[2]), .Z(n13632));
    L6MUX21 i5759 (.D0(n14293), .D1(n14294), .SD(r_addr[2]), .Z(n14301));
    L6MUX21 i5760 (.D0(n14295), .D1(n14296), .SD(r_addr[2]), .Z(n14302));
    L6MUX21 i5761 (.D0(n14297), .D1(n14298), .SD(r_addr[2]), .Z(n14303));
    L6MUX21 i5762 (.D0(n14299), .D1(n14300), .SD(r_addr[2]), .Z(n14304));
    L6MUX21 i6334 (.D0(n14871), .D1(n14872), .SD(r_addr[2]), .Z(n14876));
    L6MUX21 i5118 (.D0(n13652), .D1(n13653), .SD(r_addr[2]), .Z(n13660));
    L6MUX21 i5119 (.D0(n13654), .D1(n13655), .SD(r_addr[2]), .Z(n13661));
    L6MUX21 i5120 (.D0(n13656), .D1(n13657), .SD(r_addr[2]), .Z(n13662));
    L6MUX21 i5121 (.D0(n13658), .D1(n13659), .SD(r_addr[2]), .Z(n13663));
    L6MUX21 i6396 (.D0(n14933), .D1(n14934), .SD(r_addr[2]), .Z(n14938));
    L6MUX21 i5156 (.D0(n13690), .D1(n13691), .SD(r_addr[2]), .Z(n13698));
    L6MUX21 i5157 (.D0(n13692), .D1(n13693), .SD(r_addr[2]), .Z(n13699));
    L6MUX21 i5790 (.D0(n14324), .D1(n14325), .SD(r_addr[2]), .Z(n14332));
    L6MUX21 i5158 (.D0(n13694), .D1(n13695), .SD(r_addr[2]), .Z(n13700));
    L6MUX21 i5159 (.D0(n13696), .D1(n13697), .SD(r_addr[2]), .Z(n13701));
    L6MUX21 i5791 (.D0(n14326), .D1(n14327), .SD(r_addr[2]), .Z(n14333));
    L6MUX21 i5792 (.D0(n14328), .D1(n14329), .SD(r_addr[2]), .Z(n14334));
    L6MUX21 i5793 (.D0(n14330), .D1(n14331), .SD(r_addr[2]), .Z(n14335));
    L6MUX21 i6107 (.D0(n14641), .D1(n14642), .SD(r_addr[2]), .Z(n14649));
    L6MUX21 i6108 (.D0(n14643), .D1(n14644), .SD(r_addr[2]), .Z(n14650));
    L6MUX21 i6109 (.D0(n14645), .D1(n14646), .SD(r_addr[2]), .Z(n14651));
    L6MUX21 i6110 (.D0(n14647), .D1(n14648), .SD(r_addr[2]), .Z(n14652));
    L6MUX21 i5187 (.D0(n13721), .D1(n13722), .SD(r_addr[2]), .Z(n13729));
    L6MUX21 i5188 (.D0(n13723), .D1(n13724), .SD(r_addr[2]), .Z(n13730));
    L6MUX21 i5189 (.D0(n13725), .D1(n13726), .SD(r_addr[2]), .Z(n13731));
    L6MUX21 i5190 (.D0(n13727), .D1(n13728), .SD(r_addr[2]), .Z(n13732));
    L6MUX21 i5218 (.D0(n13752), .D1(n13753), .SD(r_addr[2]), .Z(n13760));
    L6MUX21 i5821 (.D0(n14355), .D1(n14356), .SD(r_addr[2]), .Z(n14363));
    L6MUX21 i5219 (.D0(n13754), .D1(n13755), .SD(r_addr[2]), .Z(n13761));
    L6MUX21 i5220 (.D0(n13756), .D1(n13757), .SD(r_addr[2]), .Z(n13762));
    L6MUX21 i5822 (.D0(n14357), .D1(n14358), .SD(r_addr[2]), .Z(n14364));
    L6MUX21 i5221 (.D0(n13758), .D1(n13759), .SD(r_addr[2]), .Z(n13763));
    L6MUX21 i5823 (.D0(n14359), .D1(n14360), .SD(r_addr[2]), .Z(n14365));
    L6MUX21 i5824 (.D0(n14361), .D1(n14362), .SD(r_addr[2]), .Z(n14366));
    L6MUX21 i6269 (.D0(n14803), .D1(n14804), .SD(r_addr[2]), .Z(n14811));
    L6MUX21 i6270 (.D0(n14805), .D1(n14806), .SD(r_addr[2]), .Z(n14812));
    L6MUX21 i5249 (.D0(n13783), .D1(n13784), .SD(r_addr[2]), .Z(n13791));
    L6MUX21 i5250 (.D0(n13785), .D1(n13786), .SD(r_addr[2]), .Z(n13792));
    L6MUX21 i5251 (.D0(n13787), .D1(n13788), .SD(r_addr[2]), .Z(n13793));
    L6MUX21 i6271 (.D0(n14807), .D1(n14808), .SD(r_addr[2]), .Z(n14813));
    L6MUX21 i5252 (.D0(n13789), .D1(n13790), .SD(r_addr[2]), .Z(n13794));
    L6MUX21 i6272 (.D0(n14809), .D1(n14810), .SD(r_addr[2]), .Z(n14814));
    L6MUX21 i5280 (.D0(n13814), .D1(n13815), .SD(r_addr[2]), .Z(n13822));
    L6MUX21 i5852 (.D0(n14386), .D1(n14387), .SD(r_addr[2]), .Z(n14394));
    L6MUX21 i5281 (.D0(n13816), .D1(n13817), .SD(r_addr[2]), .Z(n13823));
    L6MUX21 i5282 (.D0(n13818), .D1(n13819), .SD(r_addr[2]), .Z(n13824));
    L6MUX21 i5853 (.D0(n14388), .D1(n14389), .SD(r_addr[2]), .Z(n14395));
    L6MUX21 i5283 (.D0(n13820), .D1(n13821), .SD(r_addr[2]), .Z(n13825));
    L6MUX21 i5854 (.D0(n14390), .D1(n14391), .SD(r_addr[2]), .Z(n14396));
    L6MUX21 i5855 (.D0(n14392), .D1(n14393), .SD(r_addr[2]), .Z(n14397));
    L6MUX21 i6138 (.D0(n14672), .D1(n14673), .SD(r_addr[2]), .Z(n14680));
    L6MUX21 i6139 (.D0(n14674), .D1(n14675), .SD(r_addr[2]), .Z(n14681));
    L6MUX21 i6140 (.D0(n14676), .D1(n14677), .SD(r_addr[2]), .Z(n14682));
    L6MUX21 i6141 (.D0(n14678), .D1(n14679), .SD(r_addr[2]), .Z(n14683));
    L6MUX21 i5311 (.D0(n13845), .D1(n13846), .SD(r_addr[2]), .Z(n13853));
    L6MUX21 i5312 (.D0(n13847), .D1(n13848), .SD(r_addr[2]), .Z(n13854));
    L6MUX21 i5313 (.D0(n13849), .D1(n13850), .SD(r_addr[2]), .Z(n13855));
    L6MUX21 i5314 (.D0(n13851), .D1(n13852), .SD(r_addr[2]), .Z(n13856));
    L6MUX21 i5342 (.D0(n13876), .D1(n13877), .SD(r_addr[2]), .Z(n13884));
    L6MUX21 i5883 (.D0(n14417), .D1(n14418), .SD(r_addr[2]), .Z(n14425));
    L6MUX21 i5343 (.D0(n13878), .D1(n13879), .SD(r_addr[2]), .Z(n13885));
    L6MUX21 i5344 (.D0(n13880), .D1(n13881), .SD(r_addr[2]), .Z(n13886));
    L6MUX21 i5884 (.D0(n14419), .D1(n14420), .SD(r_addr[2]), .Z(n14426));
    L6MUX21 i5345 (.D0(n13882), .D1(n13883), .SD(r_addr[2]), .Z(n13887));
    L6MUX21 i5885 (.D0(n14421), .D1(n14422), .SD(r_addr[2]), .Z(n14427));
    L6MUX21 i5886 (.D0(n14423), .D1(n14424), .SD(r_addr[2]), .Z(n14428));
    PFUMX i4383 (.BLUT(n12909), .ALUT(n12910), .C0(r_addr[1]), .Z(n12925));
    PFUMX i4384 (.BLUT(n12911), .ALUT(n12912), .C0(r_addr[1]), .Z(n12926));
    PFUMX i4385 (.BLUT(n12913), .ALUT(n12914), .C0(r_addr[1]), .Z(n12927));
    PFUMX i4386 (.BLUT(n12915), .ALUT(n12916), .C0(r_addr[1]), .Z(n12928));
    PFUMX i4387 (.BLUT(n12917), .ALUT(n12918), .C0(r_addr[1]), .Z(n12929));
    PFUMX i5365 (.BLUT(n13891), .ALUT(n13892), .C0(r_addr[1]), .Z(n13907));
    PFUMX i4388 (.BLUT(n12919), .ALUT(n12920), .C0(r_addr[1]), .Z(n12930));
    PFUMX i4389 (.BLUT(n12921), .ALUT(n12922), .C0(r_addr[1]), .Z(n12931));
    PFUMX i5366 (.BLUT(n13893), .ALUT(n13894), .C0(r_addr[1]), .Z(n13908));
    PFUMX i4390 (.BLUT(n12923), .ALUT(n12924), .C0(r_addr[1]), .Z(n12932));
    PFUMX i5367 (.BLUT(n13895), .ALUT(n13896), .C0(r_addr[1]), .Z(n13909));
    PFUMX i5368 (.BLUT(n13897), .ALUT(n13898), .C0(r_addr[1]), .Z(n13910));
    PFUMX i5369 (.BLUT(n13899), .ALUT(n13900), .C0(r_addr[1]), .Z(n13911));
    PFUMX i5370 (.BLUT(n13901), .ALUT(n13902), .C0(r_addr[1]), .Z(n13912));
    PFUMX i5371 (.BLUT(n13903), .ALUT(n13904), .C0(r_addr[1]), .Z(n13913));
    PFUMX i5372 (.BLUT(n13905), .ALUT(n13906), .C0(r_addr[1]), .Z(n13914));
    PFUMX i4414 (.BLUT(n12940), .ALUT(n12941), .C0(r_addr[1]), .Z(n12956));
    PFUMX i4415 (.BLUT(n12942), .ALUT(n12943), .C0(r_addr[1]), .Z(n12957));
    PFUMX i4416 (.BLUT(n12944), .ALUT(n12945), .C0(r_addr[1]), .Z(n12958));
    PFUMX i4417 (.BLUT(n12946), .ALUT(n12947), .C0(r_addr[1]), .Z(n12959));
    PFUMX i4418 (.BLUT(n12948), .ALUT(n12949), .C0(r_addr[1]), .Z(n12960));
    PFUMX i4419 (.BLUT(n12950), .ALUT(n12951), .C0(r_addr[1]), .Z(n12961));
    PFUMX i4420 (.BLUT(n12952), .ALUT(n12953), .C0(r_addr[1]), .Z(n12962));
    PFUMX i4421 (.BLUT(n12954), .ALUT(n12955), .C0(r_addr[1]), .Z(n12963));
    PFUMX i4445 (.BLUT(n12971), .ALUT(n12972), .C0(r_addr[1]), .Z(n12987));
    PFUMX i4446 (.BLUT(n12973), .ALUT(n12974), .C0(r_addr[1]), .Z(n12988));
    PFUMX i4447 (.BLUT(n12975), .ALUT(n12976), .C0(r_addr[1]), .Z(n12989));
    PFUMX i4448 (.BLUT(n12977), .ALUT(n12978), .C0(r_addr[1]), .Z(n12990));
    PFUMX i4449 (.BLUT(n12979), .ALUT(n12980), .C0(r_addr[1]), .Z(n12991));
    PFUMX i4450 (.BLUT(n12981), .ALUT(n12982), .C0(r_addr[1]), .Z(n12992));
    PFUMX i4451 (.BLUT(n12983), .ALUT(n12984), .C0(r_addr[1]), .Z(n12993));
    PFUMX i4452 (.BLUT(n12985), .ALUT(n12986), .C0(r_addr[1]), .Z(n12994));
    PFUMX i5403 (.BLUT(n13929), .ALUT(n13930), .C0(r_addr[1]), .Z(n13945));
    PFUMX i5404 (.BLUT(n13931), .ALUT(n13932), .C0(r_addr[1]), .Z(n13946));
    PFUMX i5405 (.BLUT(n13933), .ALUT(n13934), .C0(r_addr[1]), .Z(n13947));
    PFUMX i5406 (.BLUT(n13935), .ALUT(n13936), .C0(r_addr[1]), .Z(n13948));
    PFUMX i5407 (.BLUT(n13937), .ALUT(n13938), .C0(r_addr[1]), .Z(n13949));
    PFUMX i5408 (.BLUT(n13939), .ALUT(n13940), .C0(r_addr[1]), .Z(n13950));
    PFUMX i4476 (.BLUT(n13002), .ALUT(n13003), .C0(r_addr[1]), .Z(n13018));
    PFUMX i5409 (.BLUT(n13941), .ALUT(n13942), .C0(r_addr[1]), .Z(n13951));
    PFUMX i4477 (.BLUT(n13004), .ALUT(n13005), .C0(r_addr[1]), .Z(n13019));
    PFUMX i4478 (.BLUT(n13006), .ALUT(n13007), .C0(r_addr[1]), .Z(n13020));
    PFUMX i5913 (.BLUT(n14439), .ALUT(n14440), .C0(r_addr[1]), .Z(n14455));
    PFUMX i5410 (.BLUT(n13943), .ALUT(n13944), .C0(r_addr[1]), .Z(n13952));
    PFUMX i4479 (.BLUT(n13008), .ALUT(n13009), .C0(r_addr[1]), .Z(n13021));
    PFUMX i4480 (.BLUT(n13010), .ALUT(n13011), .C0(r_addr[1]), .Z(n13022));
    PFUMX i4481 (.BLUT(n13012), .ALUT(n13013), .C0(r_addr[1]), .Z(n13023));
    PFUMX i4482 (.BLUT(n13014), .ALUT(n13015), .C0(r_addr[1]), .Z(n13024));
    PFUMX i5914 (.BLUT(n14441), .ALUT(n14442), .C0(r_addr[1]), .Z(n14456));
    PFUMX i4483 (.BLUT(n13016), .ALUT(n13017), .C0(r_addr[1]), .Z(n13025));
    PFUMX i5915 (.BLUT(n14443), .ALUT(n14444), .C0(r_addr[1]), .Z(n14457));
    PFUMX i5916 (.BLUT(n14445), .ALUT(n14446), .C0(r_addr[1]), .Z(n14458));
    PFUMX i5917 (.BLUT(n14447), .ALUT(n14448), .C0(r_addr[1]), .Z(n14459));
    PFUMX i5918 (.BLUT(n14449), .ALUT(n14450), .C0(r_addr[1]), .Z(n14460));
    PFUMX i5919 (.BLUT(n14451), .ALUT(n14452), .C0(r_addr[1]), .Z(n14461));
    PFUMX i6385 (.BLUT(n14911), .ALUT(n14912), .C0(r_addr[1]), .Z(n14927));
    PFUMX i6354 (.BLUT(n14880), .ALUT(n14881), .C0(r_addr[1]), .Z(n14896));
    PFUMX i6292 (.BLUT(n14818), .ALUT(n14819), .C0(r_addr[1]), .Z(n14834));
    PFUMX i6168 (.BLUT(n14694), .ALUT(n14695), .C0(r_addr[1]), .Z(n14710));
    PFUMX i5920 (.BLUT(n14453), .ALUT(n14454), .C0(r_addr[1]), .Z(n14462));
    PFUMX i4507 (.BLUT(n13033), .ALUT(n13034), .C0(r_addr[1]), .Z(n13049));
    PFUMX i4508 (.BLUT(n13035), .ALUT(n13036), .C0(r_addr[1]), .Z(n13050));
    PFUMX i4509 (.BLUT(n13037), .ALUT(n13038), .C0(r_addr[1]), .Z(n13051));
    PFUMX i4510 (.BLUT(n13039), .ALUT(n13040), .C0(r_addr[1]), .Z(n13052));
    PFUMX i4511 (.BLUT(n13041), .ALUT(n13042), .C0(r_addr[1]), .Z(n13053));
    PFUMX i4512 (.BLUT(n13043), .ALUT(n13044), .C0(r_addr[1]), .Z(n13054));
    PFUMX i4513 (.BLUT(n13045), .ALUT(n13046), .C0(r_addr[1]), .Z(n13055));
    PFUMX i4514 (.BLUT(n13047), .ALUT(n13048), .C0(r_addr[1]), .Z(n13056));
    PFUMX i6169 (.BLUT(n14696), .ALUT(n14697), .C0(r_addr[1]), .Z(n14711));
    PFUMX i6293 (.BLUT(n14820), .ALUT(n14821), .C0(r_addr[1]), .Z(n14835));
    PFUMX i6170 (.BLUT(n14698), .ALUT(n14699), .C0(r_addr[1]), .Z(n14712));
    PFUMX i5434 (.BLUT(n13960), .ALUT(n13961), .C0(r_addr[1]), .Z(n13976));
    PFUMX i5435 (.BLUT(n13962), .ALUT(n13963), .C0(r_addr[1]), .Z(n13977));
    PFUMX i5436 (.BLUT(n13964), .ALUT(n13965), .C0(r_addr[1]), .Z(n13978));
    PFUMX i6171 (.BLUT(n14700), .ALUT(n14701), .C0(r_addr[1]), .Z(n14713));
    PFUMX i5437 (.BLUT(n13966), .ALUT(n13967), .C0(r_addr[1]), .Z(n13979));
    PFUMX i5438 (.BLUT(n13968), .ALUT(n13969), .C0(r_addr[1]), .Z(n13980));
    PFUMX i5439 (.BLUT(n13970), .ALUT(n13971), .C0(r_addr[1]), .Z(n13981));
    PFUMX i5440 (.BLUT(n13972), .ALUT(n13973), .C0(r_addr[1]), .Z(n13982));
    PFUMX i6355 (.BLUT(n14882), .ALUT(n14883), .C0(r_addr[1]), .Z(n14897));
    PFUMX i6294 (.BLUT(n14822), .ALUT(n14823), .C0(r_addr[1]), .Z(n14836));
    PFUMX i6172 (.BLUT(n14702), .ALUT(n14703), .C0(r_addr[1]), .Z(n14714));
    PFUMX i5441 (.BLUT(n13974), .ALUT(n13975), .C0(r_addr[1]), .Z(n13983));
    PFUMX i6173 (.BLUT(n14704), .ALUT(n14705), .C0(r_addr[1]), .Z(n14715));
    PFUMX i6295 (.BLUT(n14824), .ALUT(n14825), .C0(r_addr[1]), .Z(n14837));
    PFUMX i6174 (.BLUT(n14706), .ALUT(n14707), .C0(r_addr[1]), .Z(n14716));
    PFUMX i6175 (.BLUT(n14708), .ALUT(n14709), .C0(r_addr[1]), .Z(n14717));
    PFUMX i6386 (.BLUT(n14913), .ALUT(n14914), .C0(r_addr[1]), .Z(n14928));
    PFUMX i6356 (.BLUT(n14884), .ALUT(n14885), .C0(r_addr[1]), .Z(n14898));
    PFUMX i6296 (.BLUT(n14826), .ALUT(n14827), .C0(r_addr[1]), .Z(n14838));
    PFUMX i5465 (.BLUT(n13991), .ALUT(n13992), .C0(r_addr[1]), .Z(n14007));
    PFUMX i6297 (.BLUT(n14828), .ALUT(n14829), .C0(r_addr[1]), .Z(n14839));
    PFUMX i5466 (.BLUT(n13993), .ALUT(n13994), .C0(r_addr[1]), .Z(n14008));
    PFUMX i5467 (.BLUT(n13995), .ALUT(n13996), .C0(r_addr[1]), .Z(n14009));
    PFUMX i5468 (.BLUT(n13997), .ALUT(n13998), .C0(r_addr[1]), .Z(n14010));
    PFUMX i5469 (.BLUT(n13999), .ALUT(n14000), .C0(r_addr[1]), .Z(n14011));
    PFUMX i5470 (.BLUT(n14001), .ALUT(n14002), .C0(r_addr[1]), .Z(n14012));
    PFUMX i5471 (.BLUT(n14003), .ALUT(n14004), .C0(r_addr[1]), .Z(n14013));
    PFUMX i5944 (.BLUT(n14470), .ALUT(n14471), .C0(r_addr[1]), .Z(n14486));
    PFUMX i5472 (.BLUT(n14005), .ALUT(n14006), .C0(r_addr[1]), .Z(n14014));
    PFUMX i6357 (.BLUT(n14886), .ALUT(n14887), .C0(r_addr[1]), .Z(n14899));
    PFUMX i6298 (.BLUT(n14830), .ALUT(n14831), .C0(r_addr[1]), .Z(n14840));
    PFUMX i5945 (.BLUT(n14472), .ALUT(n14473), .C0(r_addr[1]), .Z(n14487));
    PFUMX i5946 (.BLUT(n14474), .ALUT(n14475), .C0(r_addr[1]), .Z(n14488));
    PFUMX i4538 (.BLUT(n13064), .ALUT(n13065), .C0(r_addr[1]), .Z(n13080));
    PFUMX i4539 (.BLUT(n13066), .ALUT(n13067), .C0(r_addr[1]), .Z(n13081));
    PFUMX i5947 (.BLUT(n14476), .ALUT(n14477), .C0(r_addr[1]), .Z(n14489));
    PFUMX i4540 (.BLUT(n13068), .ALUT(n13069), .C0(r_addr[1]), .Z(n13082));
    PFUMX i4541 (.BLUT(n13070), .ALUT(n13071), .C0(r_addr[1]), .Z(n13083));
    PFUMX i4542 (.BLUT(n13072), .ALUT(n13073), .C0(r_addr[1]), .Z(n13084));
    PFUMX i4543 (.BLUT(n13074), .ALUT(n13075), .C0(r_addr[1]), .Z(n13085));
    PFUMX i5948 (.BLUT(n14478), .ALUT(n14479), .C0(r_addr[1]), .Z(n14490));
    PFUMX i4544 (.BLUT(n13076), .ALUT(n13077), .C0(r_addr[1]), .Z(n13086));
    PFUMX i4545 (.BLUT(n13078), .ALUT(n13079), .C0(r_addr[1]), .Z(n13087));
    PFUMX i6299 (.BLUT(n14832), .ALUT(n14833), .C0(r_addr[1]), .Z(n14841));
    PFUMX i5949 (.BLUT(n14480), .ALUT(n14481), .C0(r_addr[1]), .Z(n14491));
    PFUMX i5950 (.BLUT(n14482), .ALUT(n14483), .C0(r_addr[1]), .Z(n14492));
    PFUMX i5951 (.BLUT(n14484), .ALUT(n14485), .C0(r_addr[1]), .Z(n14493));
    PFUMX i6387 (.BLUT(n14915), .ALUT(n14916), .C0(r_addr[1]), .Z(n14929));
    PFUMX i6358 (.BLUT(n14888), .ALUT(n14889), .C0(r_addr[1]), .Z(n14900));
    PFUMX i4569 (.BLUT(n13095), .ALUT(n13096), .C0(r_addr[1]), .Z(n13111));
    PFUMX i4570 (.BLUT(n13097), .ALUT(n13098), .C0(r_addr[1]), .Z(n13112));
    PFUMX i4571 (.BLUT(n13099), .ALUT(n13100), .C0(r_addr[1]), .Z(n13113));
    PFUMX i4572 (.BLUT(n13101), .ALUT(n13102), .C0(r_addr[1]), .Z(n13114));
    PFUMX i4573 (.BLUT(n13103), .ALUT(n13104), .C0(r_addr[1]), .Z(n13115));
    PFUMX i5496 (.BLUT(n14022), .ALUT(n14023), .C0(r_addr[1]), .Z(n14038));
    PFUMX i4574 (.BLUT(n13105), .ALUT(n13106), .C0(r_addr[1]), .Z(n13116));
    PFUMX i4575 (.BLUT(n13107), .ALUT(n13108), .C0(r_addr[1]), .Z(n13117));
    PFUMX i5497 (.BLUT(n14024), .ALUT(n14025), .C0(r_addr[1]), .Z(n14039));
    PFUMX i4576 (.BLUT(n13109), .ALUT(n13110), .C0(r_addr[1]), .Z(n13118));
    PFUMX i5498 (.BLUT(n14026), .ALUT(n14027), .C0(r_addr[1]), .Z(n14040));
    PFUMX i5499 (.BLUT(n14028), .ALUT(n14029), .C0(r_addr[1]), .Z(n14041));
    PFUMX i5500 (.BLUT(n14030), .ALUT(n14031), .C0(r_addr[1]), .Z(n14042));
    PFUMX i5501 (.BLUT(n14032), .ALUT(n14033), .C0(r_addr[1]), .Z(n14043));
    PFUMX i5502 (.BLUT(n14034), .ALUT(n14035), .C0(r_addr[1]), .Z(n14044));
    PFUMX i5503 (.BLUT(n14036), .ALUT(n14037), .C0(r_addr[1]), .Z(n14045));
    PFUMX i6359 (.BLUT(n14890), .ALUT(n14891), .C0(r_addr[1]), .Z(n14901));
    PFUMX i4600 (.BLUT(n13126), .ALUT(n13127), .C0(r_addr[1]), .Z(n13142));
    PFUMX i4601 (.BLUT(n13128), .ALUT(n13129), .C0(r_addr[1]), .Z(n13143));
    PFUMX i4602 (.BLUT(n13130), .ALUT(n13131), .C0(r_addr[1]), .Z(n13144));
    PFUMX i4603 (.BLUT(n13132), .ALUT(n13133), .C0(r_addr[1]), .Z(n13145));
    PFUMX i4604 (.BLUT(n13134), .ALUT(n13135), .C0(r_addr[1]), .Z(n13146));
    PFUMX i4605 (.BLUT(n13136), .ALUT(n13137), .C0(r_addr[1]), .Z(n13147));
    PFUMX i4606 (.BLUT(n13138), .ALUT(n13139), .C0(r_addr[1]), .Z(n13148));
    PFUMX i4607 (.BLUT(n13140), .ALUT(n13141), .C0(r_addr[1]), .Z(n13149));
    PFUMX i6388 (.BLUT(n14917), .ALUT(n14918), .C0(r_addr[1]), .Z(n14930));
    PFUMX i6360 (.BLUT(n14892), .ALUT(n14893), .C0(r_addr[1]), .Z(n14902));
    PFUMX i5527 (.BLUT(n14053), .ALUT(n14054), .C0(r_addr[1]), .Z(n14069));
    PFUMX i5528 (.BLUT(n14055), .ALUT(n14056), .C0(r_addr[1]), .Z(n14070));
    PFUMX i4638 (.BLUT(n13164), .ALUT(n13165), .C0(r_addr[1]), .Z(n13180));
    PFUMX i4639 (.BLUT(n13166), .ALUT(n13167), .C0(r_addr[1]), .Z(n13181));
    PFUMX i5529 (.BLUT(n14057), .ALUT(n14058), .C0(r_addr[1]), .Z(n14071));
    PFUMX i4640 (.BLUT(n13168), .ALUT(n13169), .C0(r_addr[1]), .Z(n13182));
    PFUMX i4641 (.BLUT(n13170), .ALUT(n13171), .C0(r_addr[1]), .Z(n13183));
    PFUMX i5530 (.BLUT(n14059), .ALUT(n14060), .C0(r_addr[1]), .Z(n14072));
    PFUMX i4642 (.BLUT(n13172), .ALUT(n13173), .C0(r_addr[1]), .Z(n13184));
    PFUMX i4643 (.BLUT(n13174), .ALUT(n13175), .C0(r_addr[1]), .Z(n13185));
    PFUMX i5531 (.BLUT(n14061), .ALUT(n14062), .C0(r_addr[1]), .Z(n14073));
    PFUMX i4644 (.BLUT(n13176), .ALUT(n13177), .C0(r_addr[1]), .Z(n13186));
    PFUMX i4645 (.BLUT(n13178), .ALUT(n13179), .C0(r_addr[1]), .Z(n13187));
    PFUMX i5532 (.BLUT(n14063), .ALUT(n14064), .C0(r_addr[1]), .Z(n14074));
    PFUMX i5533 (.BLUT(n14065), .ALUT(n14066), .C0(r_addr[1]), .Z(n14075));
    PFUMX i5975 (.BLUT(n14501), .ALUT(n14502), .C0(r_addr[1]), .Z(n14517));
    PFUMX i5534 (.BLUT(n14067), .ALUT(n14068), .C0(r_addr[1]), .Z(n14076));
    PFUMX i5976 (.BLUT(n14503), .ALUT(n14504), .C0(r_addr[1]), .Z(n14518));
    PFUMX i5977 (.BLUT(n14505), .ALUT(n14506), .C0(r_addr[1]), .Z(n14519));
    PFUMX i6361 (.BLUT(n14894), .ALUT(n14895), .C0(r_addr[1]), .Z(n14903));
    PFUMX i5978 (.BLUT(n14507), .ALUT(n14508), .C0(r_addr[1]), .Z(n14520));
    PFUMX i5979 (.BLUT(n14509), .ALUT(n14510), .C0(r_addr[1]), .Z(n14521));
    PFUMX i4669 (.BLUT(n13195), .ALUT(n13196), .C0(r_addr[1]), .Z(n13211));
    PFUMX i4670 (.BLUT(n13197), .ALUT(n13198), .C0(r_addr[1]), .Z(n13212));
    PFUMX i5980 (.BLUT(n14511), .ALUT(n14512), .C0(r_addr[1]), .Z(n14522));
    PFUMX i4671 (.BLUT(n13199), .ALUT(n13200), .C0(r_addr[1]), .Z(n13213));
    PFUMX i4672 (.BLUT(n13201), .ALUT(n13202), .C0(r_addr[1]), .Z(n13214));
    PFUMX i4673 (.BLUT(n13203), .ALUT(n13204), .C0(r_addr[1]), .Z(n13215));
    PFUMX i4674 (.BLUT(n13205), .ALUT(n13206), .C0(r_addr[1]), .Z(n13216));
    PFUMX i5981 (.BLUT(n14513), .ALUT(n14514), .C0(r_addr[1]), .Z(n14523));
    PFUMX i4675 (.BLUT(n13207), .ALUT(n13208), .C0(r_addr[1]), .Z(n13217));
    PFUMX i4676 (.BLUT(n13209), .ALUT(n13210), .C0(r_addr[1]), .Z(n13218));
    PFUMX i6199 (.BLUT(n14725), .ALUT(n14726), .C0(r_addr[1]), .Z(n14741));
    PFUMX i5982 (.BLUT(n14515), .ALUT(n14516), .C0(r_addr[1]), .Z(n14524));
    PFUMX i6200 (.BLUT(n14727), .ALUT(n14728), .C0(r_addr[1]), .Z(n14742));
    PFUMX i6389 (.BLUT(n14919), .ALUT(n14920), .C0(r_addr[1]), .Z(n14931));
    PFUMX i6201 (.BLUT(n14729), .ALUT(n14730), .C0(r_addr[1]), .Z(n14743));
    PFUMX i5558 (.BLUT(n14084), .ALUT(n14085), .C0(r_addr[1]), .Z(n14100));
    PFUMX i5559 (.BLUT(n14086), .ALUT(n14087), .C0(r_addr[1]), .Z(n14101));
    PFUMX i4700 (.BLUT(n13226), .ALUT(n13227), .C0(r_addr[1]), .Z(n13242));
    PFUMX i5560 (.BLUT(n14088), .ALUT(n14089), .C0(r_addr[1]), .Z(n14102));
    PFUMX i4701 (.BLUT(n13228), .ALUT(n13229), .C0(r_addr[1]), .Z(n13243));
    PFUMX i4702 (.BLUT(n13230), .ALUT(n13231), .C0(r_addr[1]), .Z(n13244));
    PFUMX i6202 (.BLUT(n14731), .ALUT(n14732), .C0(r_addr[1]), .Z(n14744));
    PFUMX i5561 (.BLUT(n14090), .ALUT(n14091), .C0(r_addr[1]), .Z(n14103));
    PFUMX i4703 (.BLUT(n13232), .ALUT(n13233), .C0(r_addr[1]), .Z(n13245));
    PFUMX i4704 (.BLUT(n13234), .ALUT(n13235), .C0(r_addr[1]), .Z(n13246));
    PFUMX i5562 (.BLUT(n14092), .ALUT(n14093), .C0(r_addr[1]), .Z(n14104));
    PFUMX i4705 (.BLUT(n13236), .ALUT(n13237), .C0(r_addr[1]), .Z(n13247));
    PFUMX i4706 (.BLUT(n13238), .ALUT(n13239), .C0(r_addr[1]), .Z(n13248));
    PFUMX i5563 (.BLUT(n14094), .ALUT(n14095), .C0(r_addr[1]), .Z(n14105));
    PFUMX i4707 (.BLUT(n13240), .ALUT(n13241), .C0(r_addr[1]), .Z(n13249));
    PFUMX i5564 (.BLUT(n14096), .ALUT(n14097), .C0(r_addr[1]), .Z(n14106));
    PFUMX i6203 (.BLUT(n14733), .ALUT(n14734), .C0(r_addr[1]), .Z(n14745));
    PFUMX i5565 (.BLUT(n14098), .ALUT(n14099), .C0(r_addr[1]), .Z(n14107));
    PFUMX i6204 (.BLUT(n14735), .ALUT(n14736), .C0(r_addr[1]), .Z(n14746));
    PFUMX i6205 (.BLUT(n14737), .ALUT(n14738), .C0(r_addr[1]), .Z(n14747));
    PFUMX i4731 (.BLUT(n13257), .ALUT(n13258), .C0(r_addr[1]), .Z(n13273));
    PFUMX i4732 (.BLUT(n13259), .ALUT(n13260), .C0(r_addr[1]), .Z(n13274));
    PFUMX i4733 (.BLUT(n13261), .ALUT(n13262), .C0(r_addr[1]), .Z(n13275));
    PFUMX i4734 (.BLUT(n13263), .ALUT(n13264), .C0(r_addr[1]), .Z(n13276));
    PFUMX i4735 (.BLUT(n13265), .ALUT(n13266), .C0(r_addr[1]), .Z(n13277));
    PFUMX i6206 (.BLUT(n14739), .ALUT(n14740), .C0(r_addr[1]), .Z(n14748));
    PFUMX i4736 (.BLUT(n13267), .ALUT(n13268), .C0(r_addr[1]), .Z(n13278));
    PFUMX i4737 (.BLUT(n13269), .ALUT(n13270), .C0(r_addr[1]), .Z(n13279));
    PFUMX i4738 (.BLUT(n13271), .ALUT(n13272), .C0(r_addr[1]), .Z(n13280));
    PFUMX i5589 (.BLUT(n14115), .ALUT(n14116), .C0(r_addr[1]), .Z(n14131));
    PFUMX i6390 (.BLUT(n14921), .ALUT(n14922), .C0(r_addr[1]), .Z(n14932));
    PFUMX i5590 (.BLUT(n14117), .ALUT(n14118), .C0(r_addr[1]), .Z(n14132));
    PFUMX i4762 (.BLUT(n13288), .ALUT(n13289), .C0(r_addr[1]), .Z(n13304));
    PFUMX i5591 (.BLUT(n14119), .ALUT(n14120), .C0(r_addr[1]), .Z(n14133));
    PFUMX i4763 (.BLUT(n13290), .ALUT(n13291), .C0(r_addr[1]), .Z(n13305));
    PFUMX i4764 (.BLUT(n13292), .ALUT(n13293), .C0(r_addr[1]), .Z(n13306));
    PFUMX i5592 (.BLUT(n14121), .ALUT(n14122), .C0(r_addr[1]), .Z(n14134));
    PFUMX i4765 (.BLUT(n13294), .ALUT(n13295), .C0(r_addr[1]), .Z(n13307));
    PFUMX i4766 (.BLUT(n13296), .ALUT(n13297), .C0(r_addr[1]), .Z(n13308));
    PFUMX i5593 (.BLUT(n14123), .ALUT(n14124), .C0(r_addr[1]), .Z(n14135));
    PFUMX i4767 (.BLUT(n13298), .ALUT(n13299), .C0(r_addr[1]), .Z(n13309));
    PFUMX i4768 (.BLUT(n13300), .ALUT(n13301), .C0(r_addr[1]), .Z(n13310));
    PFUMX i5594 (.BLUT(n14125), .ALUT(n14126), .C0(r_addr[1]), .Z(n14136));
    PFUMX i4769 (.BLUT(n13302), .ALUT(n13303), .C0(r_addr[1]), .Z(n13311));
    PFUMX i5595 (.BLUT(n14127), .ALUT(n14128), .C0(r_addr[1]), .Z(n14137));
    PFUMX i6006 (.BLUT(n14532), .ALUT(n14533), .C0(r_addr[1]), .Z(n14548));
    PFUMX i5596 (.BLUT(n14129), .ALUT(n14130), .C0(r_addr[1]), .Z(n14138));
    PFUMX i6007 (.BLUT(n14534), .ALUT(n14535), .C0(r_addr[1]), .Z(n14549));
    PFUMX i6008 (.BLUT(n14536), .ALUT(n14537), .C0(r_addr[1]), .Z(n14550));
    PFUMX i6009 (.BLUT(n14538), .ALUT(n14539), .C0(r_addr[1]), .Z(n14551));
    PFUMX i6010 (.BLUT(n14540), .ALUT(n14541), .C0(r_addr[1]), .Z(n14552));
    PFUMX i4793 (.BLUT(n13319), .ALUT(n13320), .C0(r_addr[1]), .Z(n13335));
    PFUMX i6011 (.BLUT(n14542), .ALUT(n14543), .C0(r_addr[1]), .Z(n14553));
    PFUMX i4794 (.BLUT(n13321), .ALUT(n13322), .C0(r_addr[1]), .Z(n13336));
    PFUMX i4795 (.BLUT(n13323), .ALUT(n13324), .C0(r_addr[1]), .Z(n13337));
    PFUMX i4796 (.BLUT(n13325), .ALUT(n13326), .C0(r_addr[1]), .Z(n13338));
    PFUMX i4797 (.BLUT(n13327), .ALUT(n13328), .C0(r_addr[1]), .Z(n13339));
    PFUMX i6012 (.BLUT(n14544), .ALUT(n14545), .C0(r_addr[1]), .Z(n14554));
    PFUMX i4798 (.BLUT(n13329), .ALUT(n13330), .C0(r_addr[1]), .Z(n13340));
    PFUMX i4799 (.BLUT(n13331), .ALUT(n13332), .C0(r_addr[1]), .Z(n13341));
    PFUMX i4800 (.BLUT(n13333), .ALUT(n13334), .C0(r_addr[1]), .Z(n13342));
    PFUMX i6013 (.BLUT(n14546), .ALUT(n14547), .C0(r_addr[1]), .Z(n14555));
    PFUMX i5620 (.BLUT(n14146), .ALUT(n14147), .C0(r_addr[1]), .Z(n14162));
    PFUMX i5621 (.BLUT(n14148), .ALUT(n14149), .C0(r_addr[1]), .Z(n14163));
    PFUMX i4824 (.BLUT(n13350), .ALUT(n13351), .C0(r_addr[1]), .Z(n13366));
    PFUMX i5622 (.BLUT(n14150), .ALUT(n14151), .C0(r_addr[1]), .Z(n14164));
    PFUMX i4825 (.BLUT(n13352), .ALUT(n13353), .C0(r_addr[1]), .Z(n13367));
    PFUMX i6391 (.BLUT(n14923), .ALUT(n14924), .C0(r_addr[1]), .Z(n14933));
    PFUMX i5623 (.BLUT(n14152), .ALUT(n14153), .C0(r_addr[1]), .Z(n14165));
    PFUMX i4826 (.BLUT(n13354), .ALUT(n13355), .C0(r_addr[1]), .Z(n13368));
    PFUMX i4827 (.BLUT(n13356), .ALUT(n13357), .C0(r_addr[1]), .Z(n13369));
    PFUMX i5624 (.BLUT(n14154), .ALUT(n14155), .C0(r_addr[1]), .Z(n14166));
    PFUMX i4828 (.BLUT(n13358), .ALUT(n13359), .C0(r_addr[1]), .Z(n13370));
    PFUMX i4829 (.BLUT(n13360), .ALUT(n13361), .C0(r_addr[1]), .Z(n13371));
    PFUMX i5625 (.BLUT(n14156), .ALUT(n14157), .C0(r_addr[1]), .Z(n14167));
    PFUMX i4830 (.BLUT(n13362), .ALUT(n13363), .C0(r_addr[1]), .Z(n13372));
    PFUMX i4831 (.BLUT(n13364), .ALUT(n13365), .C0(r_addr[1]), .Z(n13373));
    PFUMX i5626 (.BLUT(n14158), .ALUT(n14159), .C0(r_addr[1]), .Z(n14168));
    PFUMX i5627 (.BLUT(n14160), .ALUT(n14161), .C0(r_addr[1]), .Z(n14169));
    PFUMX i4855 (.BLUT(n13381), .ALUT(n13382), .C0(r_addr[1]), .Z(n13397));
    PFUMX i4856 (.BLUT(n13383), .ALUT(n13384), .C0(r_addr[1]), .Z(n13398));
    PFUMX i4857 (.BLUT(n13385), .ALUT(n13386), .C0(r_addr[1]), .Z(n13399));
    PFUMX i4858 (.BLUT(n13387), .ALUT(n13388), .C0(r_addr[1]), .Z(n13400));
    PFUMX i4859 (.BLUT(n13389), .ALUT(n13390), .C0(r_addr[1]), .Z(n13401));
    PFUMX i4860 (.BLUT(n13391), .ALUT(n13392), .C0(r_addr[1]), .Z(n13402));
    PFUMX i4861 (.BLUT(n13393), .ALUT(n13394), .C0(r_addr[1]), .Z(n13403));
    PFUMX i4862 (.BLUT(n13395), .ALUT(n13396), .C0(r_addr[1]), .Z(n13404));
    PFUMX i6392 (.BLUT(n14925), .ALUT(n14926), .C0(r_addr[1]), .Z(n14934));
    PFUMX i4893 (.BLUT(n13419), .ALUT(n13420), .C0(r_addr[1]), .Z(n13435));
    PFUMX i4894 (.BLUT(n13421), .ALUT(n13422), .C0(r_addr[1]), .Z(n13436));
    PFUMX i4895 (.BLUT(n13423), .ALUT(n13424), .C0(r_addr[1]), .Z(n13437));
    PFUMX i6037 (.BLUT(n14563), .ALUT(n14564), .C0(r_addr[1]), .Z(n14579));
    PFUMX i5658 (.BLUT(n14184), .ALUT(n14185), .C0(r_addr[1]), .Z(n14200));
    PFUMX i4896 (.BLUT(n13425), .ALUT(n13426), .C0(r_addr[1]), .Z(n13438));
    PFUMX i4897 (.BLUT(n13427), .ALUT(n13428), .C0(r_addr[1]), .Z(n13439));
    PFUMX i5659 (.BLUT(n14186), .ALUT(n14187), .C0(r_addr[1]), .Z(n14201));
    PFUMX i4898 (.BLUT(n13429), .ALUT(n13430), .C0(r_addr[1]), .Z(n13440));
    PFUMX i4899 (.BLUT(n13431), .ALUT(n13432), .C0(r_addr[1]), .Z(n13441));
    PFUMX i6038 (.BLUT(n14565), .ALUT(n14566), .C0(r_addr[1]), .Z(n14580));
    PFUMX i5660 (.BLUT(n14188), .ALUT(n14189), .C0(r_addr[1]), .Z(n14202));
    PFUMX i4900 (.BLUT(n13433), .ALUT(n13434), .C0(r_addr[1]), .Z(n13442));
    PFUMX i5661 (.BLUT(n14190), .ALUT(n14191), .C0(r_addr[1]), .Z(n14203));
    PFUMX i6039 (.BLUT(n14567), .ALUT(n14568), .C0(r_addr[1]), .Z(n14581));
    PFUMX i5662 (.BLUT(n14192), .ALUT(n14193), .C0(r_addr[1]), .Z(n14204));
    PFUMX i5663 (.BLUT(n14194), .ALUT(n14195), .C0(r_addr[1]), .Z(n14205));
    PFUMX i6040 (.BLUT(n14569), .ALUT(n14570), .C0(r_addr[1]), .Z(n14582));
    PFUMX i5664 (.BLUT(n14196), .ALUT(n14197), .C0(r_addr[1]), .Z(n14206));
    PFUMX i5665 (.BLUT(n14198), .ALUT(n14199), .C0(r_addr[1]), .Z(n14207));
    PFUMX i6041 (.BLUT(n14571), .ALUT(n14572), .C0(r_addr[1]), .Z(n14583));
    PFUMX i6042 (.BLUT(n14573), .ALUT(n14574), .C0(r_addr[1]), .Z(n14584));
    PFUMX i6043 (.BLUT(n14575), .ALUT(n14576), .C0(r_addr[1]), .Z(n14585));
    PFUMX i4924 (.BLUT(n13450), .ALUT(n13451), .C0(r_addr[1]), .Z(n13466));
    PFUMX i6323 (.BLUT(n14849), .ALUT(n14850), .C0(r_addr[1]), .Z(n14865));
    PFUMX i6230 (.BLUT(n14756), .ALUT(n14757), .C0(r_addr[1]), .Z(n14772));
    PFUMX i6044 (.BLUT(n14577), .ALUT(n14578), .C0(r_addr[1]), .Z(n14586));
    PFUMX i4925 (.BLUT(n13452), .ALUT(n13453), .C0(r_addr[1]), .Z(n13467));
    PFUMX i4926 (.BLUT(n13454), .ALUT(n13455), .C0(r_addr[1]), .Z(n13468));
    PFUMX i4927 (.BLUT(n13456), .ALUT(n13457), .C0(r_addr[1]), .Z(n13469));
    PFUMX i4928 (.BLUT(n13458), .ALUT(n13459), .C0(r_addr[1]), .Z(n13470));
    PFUMX i4929 (.BLUT(n13460), .ALUT(n13461), .C0(r_addr[1]), .Z(n13471));
    PFUMX i4930 (.BLUT(n13462), .ALUT(n13463), .C0(r_addr[1]), .Z(n13472));
    PFUMX i4931 (.BLUT(n13464), .ALUT(n13465), .C0(r_addr[1]), .Z(n13473));
    PFUMX i6231 (.BLUT(n14758), .ALUT(n14759), .C0(r_addr[1]), .Z(n14773));
    PFUMX i6324 (.BLUT(n14851), .ALUT(n14852), .C0(r_addr[1]), .Z(n14866));
    PFUMX i6232 (.BLUT(n14760), .ALUT(n14761), .C0(r_addr[1]), .Z(n14774));
    PFUMX i6233 (.BLUT(n14762), .ALUT(n14763), .C0(r_addr[1]), .Z(n14775));
    PFUMX i4955 (.BLUT(n13481), .ALUT(n13482), .C0(r_addr[1]), .Z(n13497));
    PFUMX i4956 (.BLUT(n13483), .ALUT(n13484), .C0(r_addr[1]), .Z(n13498));
    PFUMX i6325 (.BLUT(n14853), .ALUT(n14854), .C0(r_addr[1]), .Z(n14867));
    PFUMX i6234 (.BLUT(n14764), .ALUT(n14765), .C0(r_addr[1]), .Z(n14776));
    PFUMX i5689 (.BLUT(n14215), .ALUT(n14216), .C0(r_addr[1]), .Z(n14231));
    PFUMX i4957 (.BLUT(n13485), .ALUT(n13486), .C0(r_addr[1]), .Z(n13499));
    PFUMX i4958 (.BLUT(n13487), .ALUT(n13488), .C0(r_addr[1]), .Z(n13500));
    PFUMX i5690 (.BLUT(n14217), .ALUT(n14218), .C0(r_addr[1]), .Z(n14232));
    PFUMX i4959 (.BLUT(n13489), .ALUT(n13490), .C0(r_addr[1]), .Z(n13501));
    PFUMX i4960 (.BLUT(n13491), .ALUT(n13492), .C0(r_addr[1]), .Z(n13502));
    PFUMX i5691 (.BLUT(n14219), .ALUT(n14220), .C0(r_addr[1]), .Z(n14233));
    PFUMX i4961 (.BLUT(n13493), .ALUT(n13494), .C0(r_addr[1]), .Z(n13503));
    PFUMX i4962 (.BLUT(n13495), .ALUT(n13496), .C0(r_addr[1]), .Z(n13504));
    PFUMX i5692 (.BLUT(n14221), .ALUT(n14222), .C0(r_addr[1]), .Z(n14234));
    PFUMX i6235 (.BLUT(n14766), .ALUT(n14767), .C0(r_addr[1]), .Z(n14777));
    PFUMX i5693 (.BLUT(n14223), .ALUT(n14224), .C0(r_addr[1]), .Z(n14235));
    PFUMX i5694 (.BLUT(n14225), .ALUT(n14226), .C0(r_addr[1]), .Z(n14236));
    PFUMX i5695 (.BLUT(n14227), .ALUT(n14228), .C0(r_addr[1]), .Z(n14237));
    PFUMX i5696 (.BLUT(n14229), .ALUT(n14230), .C0(r_addr[1]), .Z(n14238));
    PFUMX i6326 (.BLUT(n14855), .ALUT(n14856), .C0(r_addr[1]), .Z(n14868));
    PFUMX i6236 (.BLUT(n14768), .ALUT(n14769), .C0(r_addr[1]), .Z(n14778));
    PFUMX i6237 (.BLUT(n14770), .ALUT(n14771), .C0(r_addr[1]), .Z(n14779));
    PFUMX i4986 (.BLUT(n13512), .ALUT(n13513), .C0(r_addr[1]), .Z(n13528));
    PFUMX i4987 (.BLUT(n13514), .ALUT(n13515), .C0(r_addr[1]), .Z(n13529));
    PFUMX i4988 (.BLUT(n13516), .ALUT(n13517), .C0(r_addr[1]), .Z(n13530));
    PFUMX i4989 (.BLUT(n13518), .ALUT(n13519), .C0(r_addr[1]), .Z(n13531));
    PFUMX i6327 (.BLUT(n14857), .ALUT(n14858), .C0(r_addr[1]), .Z(n14869));
    PFUMX i4990 (.BLUT(n13520), .ALUT(n13521), .C0(r_addr[1]), .Z(n13532));
    PFUMX i4991 (.BLUT(n13522), .ALUT(n13523), .C0(r_addr[1]), .Z(n13533));
    PFUMX i4992 (.BLUT(n13524), .ALUT(n13525), .C0(r_addr[1]), .Z(n13534));
    PFUMX i4993 (.BLUT(n13526), .ALUT(n13527), .C0(r_addr[1]), .Z(n13535));
    PFUMX i6328 (.BLUT(n14859), .ALUT(n14860), .C0(r_addr[1]), .Z(n14870));
    PFUMX i5017 (.BLUT(n13543), .ALUT(n13544), .C0(r_addr[1]), .Z(n13559));
    PFUMX i5018 (.BLUT(n13545), .ALUT(n13546), .C0(r_addr[1]), .Z(n13560));
    PFUMX i6068 (.BLUT(n14594), .ALUT(n14595), .C0(r_addr[1]), .Z(n14610));
    PFUMX i5720 (.BLUT(n14246), .ALUT(n14247), .C0(r_addr[1]), .Z(n14262));
    PFUMX i5019 (.BLUT(n13547), .ALUT(n13548), .C0(r_addr[1]), .Z(n13561));
    PFUMX i5020 (.BLUT(n13549), .ALUT(n13550), .C0(r_addr[1]), .Z(n13562));
    PFUMX i5721 (.BLUT(n14248), .ALUT(n14249), .C0(r_addr[1]), .Z(n14263));
    PFUMX i5021 (.BLUT(n13551), .ALUT(n13552), .C0(r_addr[1]), .Z(n13563));
    PFUMX i5022 (.BLUT(n13553), .ALUT(n13554), .C0(r_addr[1]), .Z(n13564));
    PFUMX i6329 (.BLUT(n14861), .ALUT(n14862), .C0(r_addr[1]), .Z(n14871));
    PFUMX i6069 (.BLUT(n14596), .ALUT(n14597), .C0(r_addr[1]), .Z(n14611));
    PFUMX i5722 (.BLUT(n14250), .ALUT(n14251), .C0(r_addr[1]), .Z(n14264));
    PFUMX i5023 (.BLUT(n13555), .ALUT(n13556), .C0(r_addr[1]), .Z(n13565));
    PFUMX i5024 (.BLUT(n13557), .ALUT(n13558), .C0(r_addr[1]), .Z(n13566));
    PFUMX i5723 (.BLUT(n14252), .ALUT(n14253), .C0(r_addr[1]), .Z(n14265));
    PFUMX i6070 (.BLUT(n14598), .ALUT(n14599), .C0(r_addr[1]), .Z(n14612));
    PFUMX i5724 (.BLUT(n14254), .ALUT(n14255), .C0(r_addr[1]), .Z(n14266));
    PFUMX i5725 (.BLUT(n14256), .ALUT(n14257), .C0(r_addr[1]), .Z(n14267));
    PFUMX i6071 (.BLUT(n14600), .ALUT(n14601), .C0(r_addr[1]), .Z(n14613));
    PFUMX i5726 (.BLUT(n14258), .ALUT(n14259), .C0(r_addr[1]), .Z(n14268));
    PFUMX i5727 (.BLUT(n14260), .ALUT(n14261), .C0(r_addr[1]), .Z(n14269));
    PFUMX i6072 (.BLUT(n14602), .ALUT(n14603), .C0(r_addr[1]), .Z(n14614));
    PFUMX i6330 (.BLUT(n14863), .ALUT(n14864), .C0(r_addr[1]), .Z(n14872));
    PFUMX i6073 (.BLUT(n14604), .ALUT(n14605), .C0(r_addr[1]), .Z(n14615));
    PFUMX i6074 (.BLUT(n14606), .ALUT(n14607), .C0(r_addr[1]), .Z(n14616));
    PFUMX i6075 (.BLUT(n14608), .ALUT(n14609), .C0(r_addr[1]), .Z(n14617));
    PFUMX i5048 (.BLUT(n13574), .ALUT(n13575), .C0(r_addr[1]), .Z(n13590));
    PFUMX i5049 (.BLUT(n13576), .ALUT(n13577), .C0(r_addr[1]), .Z(n13591));
    PFUMX i5050 (.BLUT(n13578), .ALUT(n13579), .C0(r_addr[1]), .Z(n13592));
    PFUMX i5051 (.BLUT(n13580), .ALUT(n13581), .C0(r_addr[1]), .Z(n13593));
    PFUMX i5052 (.BLUT(n13582), .ALUT(n13583), .C0(r_addr[1]), .Z(n13594));
    PFUMX i5053 (.BLUT(n13584), .ALUT(n13585), .C0(r_addr[1]), .Z(n13595));
    PFUMX i5054 (.BLUT(n13586), .ALUT(n13587), .C0(r_addr[1]), .Z(n13596));
    PFUMX i5055 (.BLUT(n13588), .ALUT(n13589), .C0(r_addr[1]), .Z(n13597));
    PFUMX i5079 (.BLUT(n13605), .ALUT(n13606), .C0(r_addr[1]), .Z(n13621));
    PFUMX i5080 (.BLUT(n13607), .ALUT(n13608), .C0(r_addr[1]), .Z(n13622));
    PFUMX i5751 (.BLUT(n14277), .ALUT(n14278), .C0(r_addr[1]), .Z(n14293));
    PFUMX i5081 (.BLUT(n13609), .ALUT(n13610), .C0(r_addr[1]), .Z(n13623));
    PFUMX i5082 (.BLUT(n13611), .ALUT(n13612), .C0(r_addr[1]), .Z(n13624));
    PFUMX i5752 (.BLUT(n14279), .ALUT(n14280), .C0(r_addr[1]), .Z(n14294));
    PFUMX i5083 (.BLUT(n13613), .ALUT(n13614), .C0(r_addr[1]), .Z(n13625));
    PFUMX i5084 (.BLUT(n13615), .ALUT(n13616), .C0(r_addr[1]), .Z(n13626));
    PFUMX i5753 (.BLUT(n14281), .ALUT(n14282), .C0(r_addr[1]), .Z(n14295));
    PFUMX i5085 (.BLUT(n13617), .ALUT(n13618), .C0(r_addr[1]), .Z(n13627));
    PFUMX i5086 (.BLUT(n13619), .ALUT(n13620), .C0(r_addr[1]), .Z(n13628));
    PFUMX i5754 (.BLUT(n14283), .ALUT(n14284), .C0(r_addr[1]), .Z(n14296));
    PFUMX i5755 (.BLUT(n14285), .ALUT(n14286), .C0(r_addr[1]), .Z(n14297));
    PFUMX i5756 (.BLUT(n14287), .ALUT(n14288), .C0(r_addr[1]), .Z(n14298));
    PFUMX i5757 (.BLUT(n14289), .ALUT(n14290), .C0(r_addr[1]), .Z(n14299));
    PFUMX i5758 (.BLUT(n14291), .ALUT(n14292), .C0(r_addr[1]), .Z(n14300));
    PFUMX i5110 (.BLUT(n13636), .ALUT(n13637), .C0(r_addr[1]), .Z(n13652));
    PFUMX i5111 (.BLUT(n13638), .ALUT(n13639), .C0(r_addr[1]), .Z(n13653));
    PFUMX i5112 (.BLUT(n13640), .ALUT(n13641), .C0(r_addr[1]), .Z(n13654));
    PFUMX i5113 (.BLUT(n13642), .ALUT(n13643), .C0(r_addr[1]), .Z(n13655));
    PFUMX i5114 (.BLUT(n13644), .ALUT(n13645), .C0(r_addr[1]), .Z(n13656));
    PFUMX i5115 (.BLUT(n13646), .ALUT(n13647), .C0(r_addr[1]), .Z(n13657));
    PFUMX i5116 (.BLUT(n13648), .ALUT(n13649), .C0(r_addr[1]), .Z(n13658));
    PFUMX i5117 (.BLUT(n13650), .ALUT(n13651), .C0(r_addr[1]), .Z(n13659));
    PFUMX i6099 (.BLUT(n14625), .ALUT(n14626), .C0(r_addr[1]), .Z(n14641));
    PFUMX i5782 (.BLUT(n14308), .ALUT(n14309), .C0(r_addr[1]), .Z(n14324));
    PFUMX i5783 (.BLUT(n14310), .ALUT(n14311), .C0(r_addr[1]), .Z(n14325));
    PFUMX i6100 (.BLUT(n14627), .ALUT(n14628), .C0(r_addr[1]), .Z(n14642));
    PFUMX i5784 (.BLUT(n14312), .ALUT(n14313), .C0(r_addr[1]), .Z(n14326));
    PFUMX i5785 (.BLUT(n14314), .ALUT(n14315), .C0(r_addr[1]), .Z(n14327));
    PFUMX i5148 (.BLUT(n13674), .ALUT(n13675), .C0(r_addr[1]), .Z(n13690));
    PFUMX i5149 (.BLUT(n13676), .ALUT(n13677), .C0(r_addr[1]), .Z(n13691));
    PFUMX i6101 (.BLUT(n14629), .ALUT(n14630), .C0(r_addr[1]), .Z(n14643));
    PFUMX i5786 (.BLUT(n14316), .ALUT(n14317), .C0(r_addr[1]), .Z(n14328));
    PFUMX i5150 (.BLUT(n13678), .ALUT(n13679), .C0(r_addr[1]), .Z(n13692));
    PFUMX i5151 (.BLUT(n13680), .ALUT(n13681), .C0(r_addr[1]), .Z(n13693));
    PFUMX i5787 (.BLUT(n14318), .ALUT(n14319), .C0(r_addr[1]), .Z(n14329));
    PFUMX i5152 (.BLUT(n13682), .ALUT(n13683), .C0(r_addr[1]), .Z(n13694));
    PFUMX i5153 (.BLUT(n13684), .ALUT(n13685), .C0(r_addr[1]), .Z(n13695));
    PFUMX i6102 (.BLUT(n14631), .ALUT(n14632), .C0(r_addr[1]), .Z(n14644));
    PFUMX i5788 (.BLUT(n14320), .ALUT(n14321), .C0(r_addr[1]), .Z(n14330));
    PFUMX i5154 (.BLUT(n13686), .ALUT(n13687), .C0(r_addr[1]), .Z(n13696));
    PFUMX i5155 (.BLUT(n13688), .ALUT(n13689), .C0(r_addr[1]), .Z(n13697));
    PFUMX i5789 (.BLUT(n14322), .ALUT(n14323), .C0(r_addr[1]), .Z(n14331));
    PFUMX i6103 (.BLUT(n14633), .ALUT(n14634), .C0(r_addr[1]), .Z(n14645));
    PFUMX i6104 (.BLUT(n14635), .ALUT(n14636), .C0(r_addr[1]), .Z(n14646));
    PFUMX i6105 (.BLUT(n14637), .ALUT(n14638), .C0(r_addr[1]), .Z(n14647));
    PFUMX i6261 (.BLUT(n14787), .ALUT(n14788), .C0(r_addr[1]), .Z(n14803));
    PFUMX i6106 (.BLUT(n14639), .ALUT(n14640), .C0(r_addr[1]), .Z(n14648));
    PFUMX i6262 (.BLUT(n14789), .ALUT(n14790), .C0(r_addr[1]), .Z(n14804));
    PFUMX i5179 (.BLUT(n13705), .ALUT(n13706), .C0(r_addr[1]), .Z(n13721));
    PFUMX i5180 (.BLUT(n13707), .ALUT(n13708), .C0(r_addr[1]), .Z(n13722));
    PFUMX i5181 (.BLUT(n13709), .ALUT(n13710), .C0(r_addr[1]), .Z(n13723));
    PFUMX i5182 (.BLUT(n13711), .ALUT(n13712), .C0(r_addr[1]), .Z(n13724));
    PFUMX i5183 (.BLUT(n13713), .ALUT(n13714), .C0(r_addr[1]), .Z(n13725));
    PFUMX i5184 (.BLUT(n13715), .ALUT(n13716), .C0(r_addr[1]), .Z(n13726));
    PFUMX i5185 (.BLUT(n13717), .ALUT(n13718), .C0(r_addr[1]), .Z(n13727));
    PFUMX i5186 (.BLUT(n13719), .ALUT(n13720), .C0(r_addr[1]), .Z(n13728));
    PFUMX i6263 (.BLUT(n14791), .ALUT(n14792), .C0(r_addr[1]), .Z(n14805));
    PFUMX i6264 (.BLUT(n14793), .ALUT(n14794), .C0(r_addr[1]), .Z(n14806));
    PFUMX i6265 (.BLUT(n14795), .ALUT(n14796), .C0(r_addr[1]), .Z(n14807));
    PFUMX i5813 (.BLUT(n14339), .ALUT(n14340), .C0(r_addr[1]), .Z(n14355));
    PFUMX i5814 (.BLUT(n14341), .ALUT(n14342), .C0(r_addr[1]), .Z(n14356));
    PFUMX i5815 (.BLUT(n14343), .ALUT(n14344), .C0(r_addr[1]), .Z(n14357));
    PFUMX i5816 (.BLUT(n14345), .ALUT(n14346), .C0(r_addr[1]), .Z(n14358));
    PFUMX i5210 (.BLUT(n13736), .ALUT(n13737), .C0(r_addr[1]), .Z(n13752));
    PFUMX i5211 (.BLUT(n13738), .ALUT(n13739), .C0(r_addr[1]), .Z(n13753));
    PFUMX i6266 (.BLUT(n14797), .ALUT(n14798), .C0(r_addr[1]), .Z(n14808));
    PFUMX i5817 (.BLUT(n14347), .ALUT(n14348), .C0(r_addr[1]), .Z(n14359));
    PFUMX i5212 (.BLUT(n13740), .ALUT(n13741), .C0(r_addr[1]), .Z(n13754));
    PFUMX i5213 (.BLUT(n13742), .ALUT(n13743), .C0(r_addr[1]), .Z(n13755));
    PFUMX i5818 (.BLUT(n14349), .ALUT(n14350), .C0(r_addr[1]), .Z(n14360));
    PFUMX i5214 (.BLUT(n13744), .ALUT(n13745), .C0(r_addr[1]), .Z(n13756));
    PFUMX i5215 (.BLUT(n13746), .ALUT(n13747), .C0(r_addr[1]), .Z(n13757));
    PFUMX i5819 (.BLUT(n14351), .ALUT(n14352), .C0(r_addr[1]), .Z(n14361));
    PFUMX i5216 (.BLUT(n13748), .ALUT(n13749), .C0(r_addr[1]), .Z(n13758));
    PFUMX i5217 (.BLUT(n13750), .ALUT(n13751), .C0(r_addr[1]), .Z(n13759));
    PFUMX i5820 (.BLUT(n14353), .ALUT(n14354), .C0(r_addr[1]), .Z(n14362));
    PFUMX i6267 (.BLUT(n14799), .ALUT(n14800), .C0(r_addr[1]), .Z(n14809));
    PFUMX i6268 (.BLUT(n14801), .ALUT(n14802), .C0(r_addr[1]), .Z(n14810));
    PFUMX i5241 (.BLUT(n13767), .ALUT(n13768), .C0(r_addr[1]), .Z(n13783));
    PFUMX i5242 (.BLUT(n13769), .ALUT(n13770), .C0(r_addr[1]), .Z(n13784));
    PFUMX i5243 (.BLUT(n13771), .ALUT(n13772), .C0(r_addr[1]), .Z(n13785));
    PFUMX i5244 (.BLUT(n13773), .ALUT(n13774), .C0(r_addr[1]), .Z(n13786));
    PFUMX i5245 (.BLUT(n13775), .ALUT(n13776), .C0(r_addr[1]), .Z(n13787));
    PFUMX i5246 (.BLUT(n13777), .ALUT(n13778), .C0(r_addr[1]), .Z(n13788));
    PFUMX i5247 (.BLUT(n13779), .ALUT(n13780), .C0(r_addr[1]), .Z(n13789));
    PFUMX i5248 (.BLUT(n13781), .ALUT(n13782), .C0(r_addr[1]), .Z(n13790));
    PFUMX i6130 (.BLUT(n14656), .ALUT(n14657), .C0(r_addr[1]), .Z(n14672));
    PFUMX i5844 (.BLUT(n14370), .ALUT(n14371), .C0(r_addr[1]), .Z(n14386));
    PFUMX i5845 (.BLUT(n14372), .ALUT(n14373), .C0(r_addr[1]), .Z(n14387));
    PFUMX i6131 (.BLUT(n14658), .ALUT(n14659), .C0(r_addr[1]), .Z(n14673));
    PFUMX i5846 (.BLUT(n14374), .ALUT(n14375), .C0(r_addr[1]), .Z(n14388));
    PFUMX i5847 (.BLUT(n14376), .ALUT(n14377), .C0(r_addr[1]), .Z(n14389));
    PFUMX i5272 (.BLUT(n13798), .ALUT(n13799), .C0(r_addr[1]), .Z(n13814));
    PFUMX i6132 (.BLUT(n14660), .ALUT(n14661), .C0(r_addr[1]), .Z(n14674));
    PFUMX i5848 (.BLUT(n14378), .ALUT(n14379), .C0(r_addr[1]), .Z(n14390));
    PFUMX i5273 (.BLUT(n13800), .ALUT(n13801), .C0(r_addr[1]), .Z(n13815));
    PFUMX i5274 (.BLUT(n13802), .ALUT(n13803), .C0(r_addr[1]), .Z(n13816));
    PFUMX i5849 (.BLUT(n14380), .ALUT(n14381), .C0(r_addr[1]), .Z(n14391));
    PFUMX i5275 (.BLUT(n13804), .ALUT(n13805), .C0(r_addr[1]), .Z(n13817));
    PFUMX i5276 (.BLUT(n13806), .ALUT(n13807), .C0(r_addr[1]), .Z(n13818));
    PFUMX i6133 (.BLUT(n14662), .ALUT(n14663), .C0(r_addr[1]), .Z(n14675));
    PFUMX i5850 (.BLUT(n14382), .ALUT(n14383), .C0(r_addr[1]), .Z(n14392));
    PFUMX i5277 (.BLUT(n13808), .ALUT(n13809), .C0(r_addr[1]), .Z(n13819));
    PFUMX i5278 (.BLUT(n13810), .ALUT(n13811), .C0(r_addr[1]), .Z(n13820));
    PFUMX i5851 (.BLUT(n14384), .ALUT(n14385), .C0(r_addr[1]), .Z(n14393));
    PFUMX i5279 (.BLUT(n13812), .ALUT(n13813), .C0(r_addr[1]), .Z(n13821));
    PFUMX i6134 (.BLUT(n14664), .ALUT(n14665), .C0(r_addr[1]), .Z(n14676));
    PFUMX i6135 (.BLUT(n14666), .ALUT(n14667), .C0(r_addr[1]), .Z(n14677));
    PFUMX i6136 (.BLUT(n14668), .ALUT(n14669), .C0(r_addr[1]), .Z(n14678));
    PFUMX i6137 (.BLUT(n14670), .ALUT(n14671), .C0(r_addr[1]), .Z(n14679));
    PFUMX i5303 (.BLUT(n13829), .ALUT(n13830), .C0(r_addr[1]), .Z(n13845));
    PFUMX i5304 (.BLUT(n13831), .ALUT(n13832), .C0(r_addr[1]), .Z(n13846));
    PFUMX i5305 (.BLUT(n13833), .ALUT(n13834), .C0(r_addr[1]), .Z(n13847));
    PFUMX i5306 (.BLUT(n13835), .ALUT(n13836), .C0(r_addr[1]), .Z(n13848));
    PFUMX i5307 (.BLUT(n13837), .ALUT(n13838), .C0(r_addr[1]), .Z(n13849));
    PFUMX i5308 (.BLUT(n13839), .ALUT(n13840), .C0(r_addr[1]), .Z(n13850));
    PFUMX i5309 (.BLUT(n13841), .ALUT(n13842), .C0(r_addr[1]), .Z(n13851));
    PFUMX i5310 (.BLUT(n13843), .ALUT(n13844), .C0(r_addr[1]), .Z(n13852));
    PFUMX i5875 (.BLUT(n14401), .ALUT(n14402), .C0(r_addr[1]), .Z(n14417));
    PFUMX i5876 (.BLUT(n14403), .ALUT(n14404), .C0(r_addr[1]), .Z(n14418));
    PFUMX i5877 (.BLUT(n14405), .ALUT(n14406), .C0(r_addr[1]), .Z(n14419));
    PFUMX i5878 (.BLUT(n14407), .ALUT(n14408), .C0(r_addr[1]), .Z(n14420));
    PFUMX i5334 (.BLUT(n13860), .ALUT(n13861), .C0(r_addr[1]), .Z(n13876));
    PFUMX i5879 (.BLUT(n14409), .ALUT(n14410), .C0(r_addr[1]), .Z(n14421));
    PFUMX i5335 (.BLUT(n13862), .ALUT(n13863), .C0(r_addr[1]), .Z(n13877));
    PFUMX i5336 (.BLUT(n13864), .ALUT(n13865), .C0(r_addr[1]), .Z(n13878));
    PFUMX i5880 (.BLUT(n14411), .ALUT(n14412), .C0(r_addr[1]), .Z(n14422));
    PFUMX i5337 (.BLUT(n13866), .ALUT(n13867), .C0(r_addr[1]), .Z(n13879));
    PFUMX i5338 (.BLUT(n13868), .ALUT(n13869), .C0(r_addr[1]), .Z(n13880));
    PFUMX i5881 (.BLUT(n14413), .ALUT(n14414), .C0(r_addr[1]), .Z(n14423));
    PFUMX i5339 (.BLUT(n13870), .ALUT(n13871), .C0(r_addr[1]), .Z(n13881));
    PFUMX i5340 (.BLUT(n13872), .ALUT(n13873), .C0(r_addr[1]), .Z(n13882));
    LUT4 mux_221_i3_3_lut_4_lut (.A(n15013), .B(n14994), .C(\array[38] [2]), 
         .D(d_in_c_2), .Z(array_0__7__N_2361[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_221_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_221_i4_3_lut_4_lut (.A(n15013), .B(n14994), .C(\array[38] [3]), 
         .D(d_in_c_3), .Z(array_0__7__N_2361[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_221_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_221_i5_3_lut_4_lut (.A(n15013), .B(n14994), .C(\array[38] [4]), 
         .D(d_in_c_4), .Z(array_0__7__N_2361[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_221_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_221_i6_3_lut_4_lut (.A(n15013), .B(n14994), .C(\array[38] [5]), 
         .D(d_in_c_5), .Z(array_0__7__N_2361[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_221_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_221_i7_3_lut_4_lut (.A(n15013), .B(n14994), .C(\array[38] [6]), 
         .D(d_in_c_6), .Z(array_0__7__N_2361[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_221_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_221_i8_3_lut_4_lut (.A(n15013), .B(n14994), .C(\array[38] [7]), 
         .D(d_in_c_7), .Z(array_0__7__N_2361[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(31[11:22])
    defparam mux_221_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_4_i1_3_lut_4_lut (.A(n15023), .B(n15022), .C(\array[255] [0]), 
         .D(d_in_c_0), .Z(array_0__7__N_4097[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_4_i1_3_lut_4_lut.init = 16'hf870;
    FD1P3AX array_255___i3 (.D(array_0__7__N_4097[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[255] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i3.GSR = "ENABLED";
    FD1P3AX array_255___i4 (.D(array_0__7__N_4097[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[255] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i4.GSR = "ENABLED";
    FD1P3AX array_255___i5 (.D(array_0__7__N_4097[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[255] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i5.GSR = "ENABLED";
    FD1P3AX array_255___i6 (.D(array_0__7__N_4097[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[255] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i6.GSR = "ENABLED";
    FD1P3AX array_255___i7 (.D(array_0__7__N_4097[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[255] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i7.GSR = "ENABLED";
    FD1P3AX array_255___i8 (.D(array_0__7__N_4097[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[255] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i8.GSR = "ENABLED";
    FD1P3AX array_255___i9 (.D(array_0__7__N_4089[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[254] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i9.GSR = "ENABLED";
    FD1P3AX array_255___i10 (.D(array_0__7__N_4089[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[254] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i10.GSR = "ENABLED";
    FD1P3AX array_255___i11 (.D(array_0__7__N_4089[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[254] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i11.GSR = "ENABLED";
    FD1P3AX array_255___i12 (.D(array_0__7__N_4089[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[254] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i12.GSR = "ENABLED";
    FD1P3AX array_255___i13 (.D(array_0__7__N_4089[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[254] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i13.GSR = "ENABLED";
    FD1P3AX array_255___i14 (.D(array_0__7__N_4089[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[254] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i14.GSR = "ENABLED";
    FD1P3AX array_255___i15 (.D(array_0__7__N_4089[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[254] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i15.GSR = "ENABLED";
    FD1P3AX array_255___i16 (.D(array_0__7__N_4089[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[254] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i16.GSR = "ENABLED";
    FD1P3AX array_255___i17 (.D(array_0__7__N_4081[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[253] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i17.GSR = "ENABLED";
    FD1P3AX array_255___i18 (.D(array_0__7__N_4081[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[253] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i18.GSR = "ENABLED";
    FD1P3AX array_255___i19 (.D(array_0__7__N_4081[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[253] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i19.GSR = "ENABLED";
    FD1P3AX array_255___i20 (.D(array_0__7__N_4081[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[253] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i20.GSR = "ENABLED";
    FD1P3AX array_255___i21 (.D(array_0__7__N_4081[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[253] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i21.GSR = "ENABLED";
    FD1P3AX array_255___i22 (.D(array_0__7__N_4081[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[253] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i22.GSR = "ENABLED";
    FD1P3AX array_255___i23 (.D(array_0__7__N_4081[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[253] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i23.GSR = "ENABLED";
    FD1P3AX array_255___i24 (.D(array_0__7__N_4081[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[253] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i24.GSR = "ENABLED";
    FD1P3AX array_255___i25 (.D(array_0__7__N_4073[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[252] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i25.GSR = "ENABLED";
    FD1P3AX array_255___i26 (.D(array_0__7__N_4073[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[252] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i26.GSR = "ENABLED";
    FD1P3AX array_255___i27 (.D(array_0__7__N_4073[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[252] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i27.GSR = "ENABLED";
    FD1P3AX array_255___i28 (.D(array_0__7__N_4073[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[252] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i28.GSR = "ENABLED";
    FD1P3AX array_255___i29 (.D(array_0__7__N_4073[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[252] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i29.GSR = "ENABLED";
    FD1P3AX array_255___i30 (.D(array_0__7__N_4073[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[252] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i30.GSR = "ENABLED";
    FD1P3AX array_255___i31 (.D(array_0__7__N_4073[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[252] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i31.GSR = "ENABLED";
    FD1P3AX array_255___i32 (.D(array_0__7__N_4073[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[252] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i32.GSR = "ENABLED";
    FD1P3AX array_255___i33 (.D(array_0__7__N_4065[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[251] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i33.GSR = "ENABLED";
    FD1P3AX array_255___i34 (.D(array_0__7__N_4065[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[251] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i34.GSR = "ENABLED";
    FD1P3AX array_255___i35 (.D(array_0__7__N_4065[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[251] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i35.GSR = "ENABLED";
    FD1P3AX array_255___i36 (.D(array_0__7__N_4065[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[251] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i36.GSR = "ENABLED";
    FD1P3AX array_255___i37 (.D(array_0__7__N_4065[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[251] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i37.GSR = "ENABLED";
    FD1P3AX array_255___i38 (.D(array_0__7__N_4065[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[251] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i38.GSR = "ENABLED";
    FD1P3AX array_255___i39 (.D(array_0__7__N_4065[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[251] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i39.GSR = "ENABLED";
    FD1P3AX array_255___i40 (.D(array_0__7__N_4065[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[251] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i40.GSR = "ENABLED";
    FD1P3AX array_255___i41 (.D(array_0__7__N_4057[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[250] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i41.GSR = "ENABLED";
    FD1P3AX array_255___i42 (.D(array_0__7__N_4057[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[250] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i42.GSR = "ENABLED";
    FD1P3AX array_255___i43 (.D(array_0__7__N_4057[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[250] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i43.GSR = "ENABLED";
    FD1P3AX array_255___i44 (.D(array_0__7__N_4057[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[250] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i44.GSR = "ENABLED";
    FD1P3AX array_255___i45 (.D(array_0__7__N_4057[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[250] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i45.GSR = "ENABLED";
    FD1P3AX array_255___i46 (.D(array_0__7__N_4057[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[250] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i46.GSR = "ENABLED";
    FD1P3AX array_255___i47 (.D(array_0__7__N_4057[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[250] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i47.GSR = "ENABLED";
    FD1P3AX array_255___i48 (.D(array_0__7__N_4057[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[250] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i48.GSR = "ENABLED";
    FD1P3AX array_255___i49 (.D(array_0__7__N_4049[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[249] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i49.GSR = "ENABLED";
    FD1P3AX array_255___i50 (.D(array_0__7__N_4049[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[249] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i50.GSR = "ENABLED";
    FD1P3AX array_255___i51 (.D(array_0__7__N_4049[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[249] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i51.GSR = "ENABLED";
    FD1P3AX array_255___i52 (.D(array_0__7__N_4049[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[249] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i52.GSR = "ENABLED";
    FD1P3AX array_255___i53 (.D(array_0__7__N_4049[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[249] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i53.GSR = "ENABLED";
    FD1P3AX array_255___i54 (.D(array_0__7__N_4049[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[249] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i54.GSR = "ENABLED";
    FD1P3AX array_255___i55 (.D(array_0__7__N_4049[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[249] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i55.GSR = "ENABLED";
    FD1P3AX array_255___i56 (.D(array_0__7__N_4049[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[249] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i56.GSR = "ENABLED";
    FD1P3AX array_255___i57 (.D(array_0__7__N_4041[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[248] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i57.GSR = "ENABLED";
    FD1P3AX array_255___i58 (.D(array_0__7__N_4041[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[248] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i58.GSR = "ENABLED";
    FD1P3AX array_255___i59 (.D(array_0__7__N_4041[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[248] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i59.GSR = "ENABLED";
    FD1P3AX array_255___i60 (.D(array_0__7__N_4041[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[248] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i60.GSR = "ENABLED";
    FD1P3AX array_255___i61 (.D(array_0__7__N_4041[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[248] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i61.GSR = "ENABLED";
    FD1P3AX array_255___i62 (.D(array_0__7__N_4041[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[248] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i62.GSR = "ENABLED";
    FD1P3AX array_255___i63 (.D(array_0__7__N_4041[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[248] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i63.GSR = "ENABLED";
    FD1P3AX array_255___i64 (.D(array_0__7__N_4041[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[248] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i64.GSR = "ENABLED";
    FD1P3AX array_255___i65 (.D(array_0__7__N_4033[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[247] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i65.GSR = "ENABLED";
    FD1P3AX array_255___i66 (.D(array_0__7__N_4033[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[247] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i66.GSR = "ENABLED";
    FD1P3AX array_255___i67 (.D(array_0__7__N_4033[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[247] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i67.GSR = "ENABLED";
    FD1P3AX array_255___i68 (.D(array_0__7__N_4033[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[247] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i68.GSR = "ENABLED";
    FD1P3AX array_255___i69 (.D(array_0__7__N_4033[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[247] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i69.GSR = "ENABLED";
    FD1P3AX array_255___i70 (.D(array_0__7__N_4033[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[247] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i70.GSR = "ENABLED";
    FD1P3AX array_255___i71 (.D(array_0__7__N_4033[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[247] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i71.GSR = "ENABLED";
    FD1P3AX array_255___i72 (.D(array_0__7__N_4033[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[247] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i72.GSR = "ENABLED";
    FD1P3AX array_255___i73 (.D(array_0__7__N_4025[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[246] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i73.GSR = "ENABLED";
    FD1P3AX array_255___i74 (.D(array_0__7__N_4025[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[246] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i74.GSR = "ENABLED";
    FD1P3AX array_255___i75 (.D(array_0__7__N_4025[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[246] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i75.GSR = "ENABLED";
    FD1P3AX array_255___i76 (.D(array_0__7__N_4025[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[246] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i76.GSR = "ENABLED";
    FD1P3AX array_255___i77 (.D(array_0__7__N_4025[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[246] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i77.GSR = "ENABLED";
    FD1P3AX array_255___i78 (.D(array_0__7__N_4025[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[246] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i78.GSR = "ENABLED";
    FD1P3AX array_255___i79 (.D(array_0__7__N_4025[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[246] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i79.GSR = "ENABLED";
    FD1P3AX array_255___i80 (.D(array_0__7__N_4025[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[246] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i80.GSR = "ENABLED";
    FD1P3AX array_255___i81 (.D(array_0__7__N_4017[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[245] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i81.GSR = "ENABLED";
    FD1P3AX array_255___i82 (.D(array_0__7__N_4017[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[245] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i82.GSR = "ENABLED";
    FD1P3AX array_255___i83 (.D(array_0__7__N_4017[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[245] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i83.GSR = "ENABLED";
    FD1P3AX array_255___i84 (.D(array_0__7__N_4017[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[245] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i84.GSR = "ENABLED";
    FD1P3AX array_255___i85 (.D(array_0__7__N_4017[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[245] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i85.GSR = "ENABLED";
    FD1P3AX array_255___i86 (.D(array_0__7__N_4017[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[245] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i86.GSR = "ENABLED";
    FD1P3AX array_255___i87 (.D(array_0__7__N_4017[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[245] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i87.GSR = "ENABLED";
    FD1P3AX array_255___i88 (.D(array_0__7__N_4017[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[245] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i88.GSR = "ENABLED";
    FD1P3AX array_255___i89 (.D(array_0__7__N_4009[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[244] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i89.GSR = "ENABLED";
    FD1P3AX array_255___i90 (.D(array_0__7__N_4009[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[244] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i90.GSR = "ENABLED";
    FD1P3AX array_255___i91 (.D(array_0__7__N_4009[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[244] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i91.GSR = "ENABLED";
    FD1P3AX array_255___i92 (.D(array_0__7__N_4009[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[244] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i92.GSR = "ENABLED";
    FD1P3AX array_255___i93 (.D(array_0__7__N_4009[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[244] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i93.GSR = "ENABLED";
    FD1P3AX array_255___i94 (.D(array_0__7__N_4009[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[244] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i94.GSR = "ENABLED";
    FD1P3AX array_255___i95 (.D(array_0__7__N_4009[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[244] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i95.GSR = "ENABLED";
    FD1P3AX array_255___i96 (.D(array_0__7__N_4009[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[244] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i96.GSR = "ENABLED";
    FD1P3AX array_255___i97 (.D(array_0__7__N_4001[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[243] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i97.GSR = "ENABLED";
    FD1P3AX array_255___i98 (.D(array_0__7__N_4001[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[243] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i98.GSR = "ENABLED";
    FD1P3AX array_255___i99 (.D(array_0__7__N_4001[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[243] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i99.GSR = "ENABLED";
    FD1P3AX array_255___i100 (.D(array_0__7__N_4001[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[243] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i100.GSR = "ENABLED";
    FD1P3AX array_255___i101 (.D(array_0__7__N_4001[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[243] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i101.GSR = "ENABLED";
    FD1P3AX array_255___i102 (.D(array_0__7__N_4001[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[243] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i102.GSR = "ENABLED";
    FD1P3AX array_255___i103 (.D(array_0__7__N_4001[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[243] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i103.GSR = "ENABLED";
    FD1P3AX array_255___i104 (.D(array_0__7__N_4001[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[243] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i104.GSR = "ENABLED";
    FD1P3AX array_255___i105 (.D(array_0__7__N_3993[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[242] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i105.GSR = "ENABLED";
    FD1P3AX array_255___i106 (.D(array_0__7__N_3993[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[242] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i106.GSR = "ENABLED";
    FD1P3AX array_255___i107 (.D(array_0__7__N_3993[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[242] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i107.GSR = "ENABLED";
    FD1P3AX array_255___i108 (.D(array_0__7__N_3993[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[242] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i108.GSR = "ENABLED";
    FD1P3AX array_255___i109 (.D(array_0__7__N_3993[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[242] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i109.GSR = "ENABLED";
    FD1P3AX array_255___i110 (.D(array_0__7__N_3993[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[242] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i110.GSR = "ENABLED";
    FD1P3AX array_255___i111 (.D(array_0__7__N_3993[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[242] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i111.GSR = "ENABLED";
    FD1P3AX array_255___i112 (.D(array_0__7__N_3993[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[242] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i112.GSR = "ENABLED";
    FD1P3AX array_255___i113 (.D(array_0__7__N_3985[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[241] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i113.GSR = "ENABLED";
    FD1P3AX array_255___i114 (.D(array_0__7__N_3985[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[241] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i114.GSR = "ENABLED";
    FD1P3AX array_255___i115 (.D(array_0__7__N_3985[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[241] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i115.GSR = "ENABLED";
    FD1P3AX array_255___i116 (.D(array_0__7__N_3985[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[241] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i116.GSR = "ENABLED";
    FD1P3AX array_255___i117 (.D(array_0__7__N_3985[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[241] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i117.GSR = "ENABLED";
    FD1P3AX array_255___i118 (.D(array_0__7__N_3985[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[241] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i118.GSR = "ENABLED";
    FD1P3AX array_255___i119 (.D(array_0__7__N_3985[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[241] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i119.GSR = "ENABLED";
    FD1P3AX array_255___i120 (.D(array_0__7__N_3985[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[241] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i120.GSR = "ENABLED";
    FD1P3AX array_255___i121 (.D(array_0__7__N_3977[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[240] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i121.GSR = "ENABLED";
    FD1P3AX array_255___i122 (.D(array_0__7__N_3977[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[240] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i122.GSR = "ENABLED";
    FD1P3AX array_255___i123 (.D(array_0__7__N_3977[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[240] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i123.GSR = "ENABLED";
    FD1P3AX array_255___i124 (.D(array_0__7__N_3977[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[240] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i124.GSR = "ENABLED";
    FD1P3AX array_255___i125 (.D(array_0__7__N_3977[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[240] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i125.GSR = "ENABLED";
    FD1P3AX array_255___i126 (.D(array_0__7__N_3977[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[240] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i126.GSR = "ENABLED";
    FD1P3AX array_255___i127 (.D(array_0__7__N_3977[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[240] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i127.GSR = "ENABLED";
    FD1P3AX array_255___i128 (.D(array_0__7__N_3977[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[240] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i128.GSR = "ENABLED";
    FD1P3AX array_255___i129 (.D(array_0__7__N_3969[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[239] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i129.GSR = "ENABLED";
    FD1P3AX array_255___i130 (.D(array_0__7__N_3969[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[239] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i130.GSR = "ENABLED";
    FD1P3AX array_255___i131 (.D(array_0__7__N_3969[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[239] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i131.GSR = "ENABLED";
    FD1P3AX array_255___i132 (.D(array_0__7__N_3969[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[239] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i132.GSR = "ENABLED";
    FD1P3AX array_255___i133 (.D(array_0__7__N_3969[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[239] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i133.GSR = "ENABLED";
    FD1P3AX array_255___i134 (.D(array_0__7__N_3969[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[239] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i134.GSR = "ENABLED";
    FD1P3AX array_255___i135 (.D(array_0__7__N_3969[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[239] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i135.GSR = "ENABLED";
    FD1P3AX array_255___i136 (.D(array_0__7__N_3969[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[239] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i136.GSR = "ENABLED";
    FD1P3AX array_255___i137 (.D(array_0__7__N_3961[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[238] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i137.GSR = "ENABLED";
    FD1P3AX array_255___i138 (.D(array_0__7__N_3961[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[238] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i138.GSR = "ENABLED";
    FD1P3AX array_255___i139 (.D(array_0__7__N_3961[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[238] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i139.GSR = "ENABLED";
    FD1P3AX array_255___i140 (.D(array_0__7__N_3961[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[238] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i140.GSR = "ENABLED";
    FD1P3AX array_255___i141 (.D(array_0__7__N_3961[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[238] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i141.GSR = "ENABLED";
    FD1P3AX array_255___i142 (.D(array_0__7__N_3961[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[238] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i142.GSR = "ENABLED";
    FD1P3AX array_255___i143 (.D(array_0__7__N_3961[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[238] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i143.GSR = "ENABLED";
    FD1P3AX array_255___i144 (.D(array_0__7__N_3961[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[238] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i144.GSR = "ENABLED";
    FD1P3AX array_255___i145 (.D(array_0__7__N_3953[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[237] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i145.GSR = "ENABLED";
    FD1P3AX array_255___i146 (.D(array_0__7__N_3953[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[237] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i146.GSR = "ENABLED";
    FD1P3AX array_255___i147 (.D(array_0__7__N_3953[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[237] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i147.GSR = "ENABLED";
    FD1P3AX array_255___i148 (.D(array_0__7__N_3953[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[237] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i148.GSR = "ENABLED";
    FD1P3AX array_255___i149 (.D(array_0__7__N_3953[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[237] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i149.GSR = "ENABLED";
    FD1P3AX array_255___i150 (.D(array_0__7__N_3953[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[237] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i150.GSR = "ENABLED";
    FD1P3AX array_255___i151 (.D(array_0__7__N_3953[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[237] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i151.GSR = "ENABLED";
    FD1P3AX array_255___i152 (.D(array_0__7__N_3953[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[237] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i152.GSR = "ENABLED";
    FD1P3AX array_255___i153 (.D(array_0__7__N_3945[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[236] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i153.GSR = "ENABLED";
    FD1P3AX array_255___i154 (.D(array_0__7__N_3945[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[236] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i154.GSR = "ENABLED";
    FD1P3AX array_255___i155 (.D(array_0__7__N_3945[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[236] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i155.GSR = "ENABLED";
    FD1P3AX array_255___i156 (.D(array_0__7__N_3945[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[236] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i156.GSR = "ENABLED";
    FD1P3AX array_255___i157 (.D(array_0__7__N_3945[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[236] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i157.GSR = "ENABLED";
    FD1P3AX array_255___i158 (.D(array_0__7__N_3945[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[236] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i158.GSR = "ENABLED";
    FD1P3AX array_255___i159 (.D(array_0__7__N_3945[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[236] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i159.GSR = "ENABLED";
    FD1P3AX array_255___i160 (.D(array_0__7__N_3945[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[236] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i160.GSR = "ENABLED";
    FD1P3AX array_255___i161 (.D(array_0__7__N_3937[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[235] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i161.GSR = "ENABLED";
    FD1P3AX array_255___i162 (.D(array_0__7__N_3937[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[235] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i162.GSR = "ENABLED";
    FD1P3AX array_255___i163 (.D(array_0__7__N_3937[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[235] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i163.GSR = "ENABLED";
    FD1P3AX array_255___i164 (.D(array_0__7__N_3937[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[235] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i164.GSR = "ENABLED";
    FD1P3AX array_255___i165 (.D(array_0__7__N_3937[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[235] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i165.GSR = "ENABLED";
    FD1P3AX array_255___i166 (.D(array_0__7__N_3937[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[235] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i166.GSR = "ENABLED";
    FD1P3AX array_255___i167 (.D(array_0__7__N_3937[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[235] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i167.GSR = "ENABLED";
    FD1P3AX array_255___i168 (.D(array_0__7__N_3937[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[235] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i168.GSR = "ENABLED";
    FD1P3AX array_255___i169 (.D(array_0__7__N_3929[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[234] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i169.GSR = "ENABLED";
    FD1P3AX array_255___i170 (.D(array_0__7__N_3929[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[234] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i170.GSR = "ENABLED";
    FD1P3AX array_255___i171 (.D(array_0__7__N_3929[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[234] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i171.GSR = "ENABLED";
    FD1P3AX array_255___i172 (.D(array_0__7__N_3929[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[234] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i172.GSR = "ENABLED";
    FD1P3AX array_255___i173 (.D(array_0__7__N_3929[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[234] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i173.GSR = "ENABLED";
    FD1P3AX array_255___i174 (.D(array_0__7__N_3929[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[234] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i174.GSR = "ENABLED";
    FD1P3AX array_255___i175 (.D(array_0__7__N_3929[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[234] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i175.GSR = "ENABLED";
    FD1P3AX array_255___i176 (.D(array_0__7__N_3929[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[234] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i176.GSR = "ENABLED";
    FD1P3AX array_255___i177 (.D(array_0__7__N_3921[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[233] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i177.GSR = "ENABLED";
    FD1P3AX array_255___i178 (.D(array_0__7__N_3921[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[233] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i178.GSR = "ENABLED";
    FD1P3AX array_255___i179 (.D(array_0__7__N_3921[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[233] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i179.GSR = "ENABLED";
    FD1P3AX array_255___i180 (.D(array_0__7__N_3921[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[233] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i180.GSR = "ENABLED";
    FD1P3AX array_255___i181 (.D(array_0__7__N_3921[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[233] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i181.GSR = "ENABLED";
    FD1P3AX array_255___i182 (.D(array_0__7__N_3921[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[233] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i182.GSR = "ENABLED";
    FD1P3AX array_255___i183 (.D(array_0__7__N_3921[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[233] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i183.GSR = "ENABLED";
    FD1P3AX array_255___i184 (.D(array_0__7__N_3921[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[233] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i184.GSR = "ENABLED";
    FD1P3AX array_255___i185 (.D(array_0__7__N_3913[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[232] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i185.GSR = "ENABLED";
    FD1P3AX array_255___i186 (.D(array_0__7__N_3913[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[232] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i186.GSR = "ENABLED";
    FD1P3AX array_255___i187 (.D(array_0__7__N_3913[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[232] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i187.GSR = "ENABLED";
    FD1P3AX array_255___i188 (.D(array_0__7__N_3913[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[232] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i188.GSR = "ENABLED";
    FD1P3AX array_255___i189 (.D(array_0__7__N_3913[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[232] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i189.GSR = "ENABLED";
    FD1P3AX array_255___i190 (.D(array_0__7__N_3913[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[232] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i190.GSR = "ENABLED";
    FD1P3AX array_255___i191 (.D(array_0__7__N_3913[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[232] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i191.GSR = "ENABLED";
    FD1P3AX array_255___i192 (.D(array_0__7__N_3913[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[232] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i192.GSR = "ENABLED";
    FD1P3AX array_255___i193 (.D(array_0__7__N_3905[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[231] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i193.GSR = "ENABLED";
    FD1P3AX array_255___i194 (.D(array_0__7__N_3905[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[231] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i194.GSR = "ENABLED";
    FD1P3AX array_255___i195 (.D(array_0__7__N_3905[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[231] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i195.GSR = "ENABLED";
    FD1P3AX array_255___i196 (.D(array_0__7__N_3905[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[231] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i196.GSR = "ENABLED";
    FD1P3AX array_255___i197 (.D(array_0__7__N_3905[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[231] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i197.GSR = "ENABLED";
    FD1P3AX array_255___i198 (.D(array_0__7__N_3905[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[231] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i198.GSR = "ENABLED";
    FD1P3AX array_255___i199 (.D(array_0__7__N_3905[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[231] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i199.GSR = "ENABLED";
    FD1P3AX array_255___i200 (.D(array_0__7__N_3905[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[231] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i200.GSR = "ENABLED";
    FD1P3AX array_255___i201 (.D(array_0__7__N_3897[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[230] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i201.GSR = "ENABLED";
    FD1P3AX array_255___i202 (.D(array_0__7__N_3897[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[230] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i202.GSR = "ENABLED";
    FD1P3AX array_255___i203 (.D(array_0__7__N_3897[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[230] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i203.GSR = "ENABLED";
    FD1P3AX array_255___i204 (.D(array_0__7__N_3897[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[230] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i204.GSR = "ENABLED";
    FD1P3AX array_255___i205 (.D(array_0__7__N_3897[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[230] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i205.GSR = "ENABLED";
    FD1P3AX array_255___i206 (.D(array_0__7__N_3897[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[230] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i206.GSR = "ENABLED";
    FD1P3AX array_255___i207 (.D(array_0__7__N_3897[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[230] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i207.GSR = "ENABLED";
    FD1P3AX array_255___i208 (.D(array_0__7__N_3897[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[230] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i208.GSR = "ENABLED";
    FD1P3AX array_255___i209 (.D(array_0__7__N_3889[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[229] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i209.GSR = "ENABLED";
    FD1P3AX array_255___i210 (.D(array_0__7__N_3889[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[229] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i210.GSR = "ENABLED";
    FD1P3AX array_255___i211 (.D(array_0__7__N_3889[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[229] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i211.GSR = "ENABLED";
    FD1P3AX array_255___i212 (.D(array_0__7__N_3889[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[229] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i212.GSR = "ENABLED";
    FD1P3AX array_255___i213 (.D(array_0__7__N_3889[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[229] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i213.GSR = "ENABLED";
    FD1P3AX array_255___i214 (.D(array_0__7__N_3889[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[229] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i214.GSR = "ENABLED";
    FD1P3AX array_255___i215 (.D(array_0__7__N_3889[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[229] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i215.GSR = "ENABLED";
    FD1P3AX array_255___i216 (.D(array_0__7__N_3889[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[229] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i216.GSR = "ENABLED";
    FD1P3AX array_255___i217 (.D(array_0__7__N_3881[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[228] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i217.GSR = "ENABLED";
    FD1P3AX array_255___i218 (.D(array_0__7__N_3881[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[228] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i218.GSR = "ENABLED";
    FD1P3AX array_255___i219 (.D(array_0__7__N_3881[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[228] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i219.GSR = "ENABLED";
    FD1P3AX array_255___i220 (.D(array_0__7__N_3881[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[228] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i220.GSR = "ENABLED";
    FD1P3AX array_255___i221 (.D(array_0__7__N_3881[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[228] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i221.GSR = "ENABLED";
    FD1P3AX array_255___i222 (.D(array_0__7__N_3881[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[228] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i222.GSR = "ENABLED";
    FD1P3AX array_255___i223 (.D(array_0__7__N_3881[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[228] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i223.GSR = "ENABLED";
    FD1P3AX array_255___i224 (.D(array_0__7__N_3881[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[228] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i224.GSR = "ENABLED";
    FD1P3AX array_255___i225 (.D(array_0__7__N_3873[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[227] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i225.GSR = "ENABLED";
    FD1P3AX array_255___i226 (.D(array_0__7__N_3873[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[227] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i226.GSR = "ENABLED";
    FD1P3AX array_255___i227 (.D(array_0__7__N_3873[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[227] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i227.GSR = "ENABLED";
    FD1P3AX array_255___i228 (.D(array_0__7__N_3873[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[227] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i228.GSR = "ENABLED";
    FD1P3AX array_255___i229 (.D(array_0__7__N_3873[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[227] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i229.GSR = "ENABLED";
    FD1P3AX array_255___i230 (.D(array_0__7__N_3873[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[227] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i230.GSR = "ENABLED";
    FD1P3AX array_255___i231 (.D(array_0__7__N_3873[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[227] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i231.GSR = "ENABLED";
    FD1P3AX array_255___i232 (.D(array_0__7__N_3873[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[227] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i232.GSR = "ENABLED";
    FD1P3AX array_255___i233 (.D(array_0__7__N_3865[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[226] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i233.GSR = "ENABLED";
    FD1P3AX array_255___i234 (.D(array_0__7__N_3865[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[226] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i234.GSR = "ENABLED";
    FD1P3AX array_255___i235 (.D(array_0__7__N_3865[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[226] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i235.GSR = "ENABLED";
    FD1P3AX array_255___i236 (.D(array_0__7__N_3865[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[226] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i236.GSR = "ENABLED";
    FD1P3AX array_255___i237 (.D(array_0__7__N_3865[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[226] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i237.GSR = "ENABLED";
    FD1P3AX array_255___i238 (.D(array_0__7__N_3865[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[226] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i238.GSR = "ENABLED";
    FD1P3AX array_255___i239 (.D(array_0__7__N_3865[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[226] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i239.GSR = "ENABLED";
    FD1P3AX array_255___i240 (.D(array_0__7__N_3865[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[226] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i240.GSR = "ENABLED";
    FD1P3AX array_255___i241 (.D(array_0__7__N_3857[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[225] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i241.GSR = "ENABLED";
    FD1P3AX array_255___i242 (.D(array_0__7__N_3857[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[225] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i242.GSR = "ENABLED";
    FD1P3AX array_255___i243 (.D(array_0__7__N_3857[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[225] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i243.GSR = "ENABLED";
    FD1P3AX array_255___i244 (.D(array_0__7__N_3857[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[225] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i244.GSR = "ENABLED";
    FD1P3AX array_255___i245 (.D(array_0__7__N_3857[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[225] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i245.GSR = "ENABLED";
    FD1P3AX array_255___i246 (.D(array_0__7__N_3857[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[225] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i246.GSR = "ENABLED";
    FD1P3AX array_255___i247 (.D(array_0__7__N_3857[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[225] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i247.GSR = "ENABLED";
    FD1P3AX array_255___i248 (.D(array_0__7__N_3857[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[225] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i248.GSR = "ENABLED";
    FD1P3AX array_255___i249 (.D(array_0__7__N_3849[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[224] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i249.GSR = "ENABLED";
    FD1P3AX array_255___i250 (.D(array_0__7__N_3849[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[224] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i250.GSR = "ENABLED";
    FD1P3AX array_255___i251 (.D(array_0__7__N_3849[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[224] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i251.GSR = "ENABLED";
    FD1P3AX array_255___i252 (.D(array_0__7__N_3849[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[224] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i252.GSR = "ENABLED";
    FD1P3AX array_255___i253 (.D(array_0__7__N_3849[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[224] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i253.GSR = "ENABLED";
    FD1P3AX array_255___i254 (.D(array_0__7__N_3849[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[224] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i254.GSR = "ENABLED";
    FD1P3AX array_255___i255 (.D(array_0__7__N_3849[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[224] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i255.GSR = "ENABLED";
    FD1P3AX array_255___i256 (.D(array_0__7__N_3849[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[224] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i256.GSR = "ENABLED";
    FD1P3AX array_255___i257 (.D(array_0__7__N_3841[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[223] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i257.GSR = "ENABLED";
    FD1P3AX array_255___i258 (.D(array_0__7__N_3841[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[223] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i258.GSR = "ENABLED";
    FD1P3AX array_255___i259 (.D(array_0__7__N_3841[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[223] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i259.GSR = "ENABLED";
    FD1P3AX array_255___i260 (.D(array_0__7__N_3841[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[223] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i260.GSR = "ENABLED";
    FD1P3AX array_255___i261 (.D(array_0__7__N_3841[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[223] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i261.GSR = "ENABLED";
    FD1P3AX array_255___i262 (.D(array_0__7__N_3841[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[223] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i262.GSR = "ENABLED";
    FD1P3AX array_255___i263 (.D(array_0__7__N_3841[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[223] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i263.GSR = "ENABLED";
    FD1P3AX array_255___i264 (.D(array_0__7__N_3841[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[223] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i264.GSR = "ENABLED";
    FD1P3AX array_255___i265 (.D(array_0__7__N_3833[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[222] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i265.GSR = "ENABLED";
    FD1P3AX array_255___i266 (.D(array_0__7__N_3833[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[222] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i266.GSR = "ENABLED";
    FD1P3AX array_255___i267 (.D(array_0__7__N_3833[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[222] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i267.GSR = "ENABLED";
    FD1P3AX array_255___i268 (.D(array_0__7__N_3833[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[222] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i268.GSR = "ENABLED";
    FD1P3AX array_255___i269 (.D(array_0__7__N_3833[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[222] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i269.GSR = "ENABLED";
    FD1P3AX array_255___i270 (.D(array_0__7__N_3833[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[222] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i270.GSR = "ENABLED";
    FD1P3AX array_255___i271 (.D(array_0__7__N_3833[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[222] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i271.GSR = "ENABLED";
    FD1P3AX array_255___i272 (.D(array_0__7__N_3833[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[222] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i272.GSR = "ENABLED";
    FD1P3AX array_255___i273 (.D(array_0__7__N_3825[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[221] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i273.GSR = "ENABLED";
    FD1P3AX array_255___i274 (.D(array_0__7__N_3825[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[221] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i274.GSR = "ENABLED";
    FD1P3AX array_255___i275 (.D(array_0__7__N_3825[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[221] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i275.GSR = "ENABLED";
    FD1P3AX array_255___i276 (.D(array_0__7__N_3825[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[221] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i276.GSR = "ENABLED";
    FD1P3AX array_255___i277 (.D(array_0__7__N_3825[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[221] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i277.GSR = "ENABLED";
    FD1P3AX array_255___i278 (.D(array_0__7__N_3825[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[221] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i278.GSR = "ENABLED";
    FD1P3AX array_255___i279 (.D(array_0__7__N_3825[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[221] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i279.GSR = "ENABLED";
    FD1P3AX array_255___i280 (.D(array_0__7__N_3825[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[221] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i280.GSR = "ENABLED";
    FD1P3AX array_255___i281 (.D(array_0__7__N_3817[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[220] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i281.GSR = "ENABLED";
    FD1P3AX array_255___i282 (.D(array_0__7__N_3817[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[220] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i282.GSR = "ENABLED";
    FD1P3AX array_255___i283 (.D(array_0__7__N_3817[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[220] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i283.GSR = "ENABLED";
    FD1P3AX array_255___i284 (.D(array_0__7__N_3817[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[220] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i284.GSR = "ENABLED";
    FD1P3AX array_255___i285 (.D(array_0__7__N_3817[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[220] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i285.GSR = "ENABLED";
    FD1P3AX array_255___i286 (.D(array_0__7__N_3817[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[220] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i286.GSR = "ENABLED";
    FD1P3AX array_255___i287 (.D(array_0__7__N_3817[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[220] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i287.GSR = "ENABLED";
    FD1P3AX array_255___i288 (.D(array_0__7__N_3817[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[220] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i288.GSR = "ENABLED";
    FD1P3AX array_255___i289 (.D(array_0__7__N_3809[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[219] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i289.GSR = "ENABLED";
    FD1P3AX array_255___i290 (.D(array_0__7__N_3809[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[219] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i290.GSR = "ENABLED";
    FD1P3AX array_255___i291 (.D(array_0__7__N_3809[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[219] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i291.GSR = "ENABLED";
    FD1P3AX array_255___i292 (.D(array_0__7__N_3809[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[219] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i292.GSR = "ENABLED";
    FD1P3AX array_255___i293 (.D(array_0__7__N_3809[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[219] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i293.GSR = "ENABLED";
    FD1P3AX array_255___i294 (.D(array_0__7__N_3809[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[219] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i294.GSR = "ENABLED";
    FD1P3AX array_255___i295 (.D(array_0__7__N_3809[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[219] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i295.GSR = "ENABLED";
    FD1P3AX array_255___i296 (.D(array_0__7__N_3809[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[219] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i296.GSR = "ENABLED";
    FD1P3AX array_255___i297 (.D(array_0__7__N_3801[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[218] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i297.GSR = "ENABLED";
    FD1P3AX array_255___i298 (.D(array_0__7__N_3801[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[218] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i298.GSR = "ENABLED";
    FD1P3AX array_255___i299 (.D(array_0__7__N_3801[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[218] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i299.GSR = "ENABLED";
    FD1P3AX array_255___i300 (.D(array_0__7__N_3801[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[218] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i300.GSR = "ENABLED";
    FD1P3AX array_255___i301 (.D(array_0__7__N_3801[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[218] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i301.GSR = "ENABLED";
    FD1P3AX array_255___i302 (.D(array_0__7__N_3801[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[218] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i302.GSR = "ENABLED";
    FD1P3AX array_255___i303 (.D(array_0__7__N_3801[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[218] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i303.GSR = "ENABLED";
    FD1P3AX array_255___i304 (.D(array_0__7__N_3801[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[218] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i304.GSR = "ENABLED";
    FD1P3AX array_255___i305 (.D(array_0__7__N_3793[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[217] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i305.GSR = "ENABLED";
    FD1P3AX array_255___i306 (.D(array_0__7__N_3793[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[217] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i306.GSR = "ENABLED";
    FD1P3AX array_255___i307 (.D(array_0__7__N_3793[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[217] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i307.GSR = "ENABLED";
    FD1P3AX array_255___i308 (.D(array_0__7__N_3793[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[217] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i308.GSR = "ENABLED";
    FD1P3AX array_255___i309 (.D(array_0__7__N_3793[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[217] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i309.GSR = "ENABLED";
    FD1P3AX array_255___i310 (.D(array_0__7__N_3793[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[217] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i310.GSR = "ENABLED";
    FD1P3AX array_255___i311 (.D(array_0__7__N_3793[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[217] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i311.GSR = "ENABLED";
    FD1P3AX array_255___i312 (.D(array_0__7__N_3793[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[217] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i312.GSR = "ENABLED";
    FD1P3AX array_255___i313 (.D(array_0__7__N_3785[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[216] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i313.GSR = "ENABLED";
    FD1P3AX array_255___i314 (.D(array_0__7__N_3785[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[216] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i314.GSR = "ENABLED";
    FD1P3AX array_255___i315 (.D(array_0__7__N_3785[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[216] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i315.GSR = "ENABLED";
    FD1P3AX array_255___i316 (.D(array_0__7__N_3785[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[216] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i316.GSR = "ENABLED";
    FD1P3AX array_255___i317 (.D(array_0__7__N_3785[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[216] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i317.GSR = "ENABLED";
    FD1P3AX array_255___i318 (.D(array_0__7__N_3785[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[216] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i318.GSR = "ENABLED";
    FD1P3AX array_255___i319 (.D(array_0__7__N_3785[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[216] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i319.GSR = "ENABLED";
    FD1P3AX array_255___i320 (.D(array_0__7__N_3785[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[216] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i320.GSR = "ENABLED";
    FD1P3AX array_255___i321 (.D(array_0__7__N_3777[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[215] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i321.GSR = "ENABLED";
    FD1P3AX array_255___i322 (.D(array_0__7__N_3777[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[215] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i322.GSR = "ENABLED";
    FD1P3AX array_255___i323 (.D(array_0__7__N_3777[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[215] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i323.GSR = "ENABLED";
    FD1P3AX array_255___i324 (.D(array_0__7__N_3777[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[215] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i324.GSR = "ENABLED";
    FD1P3AX array_255___i325 (.D(array_0__7__N_3777[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[215] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i325.GSR = "ENABLED";
    FD1P3AX array_255___i326 (.D(array_0__7__N_3777[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[215] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i326.GSR = "ENABLED";
    FD1P3AX array_255___i327 (.D(array_0__7__N_3777[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[215] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i327.GSR = "ENABLED";
    FD1P3AX array_255___i328 (.D(array_0__7__N_3777[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[215] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i328.GSR = "ENABLED";
    FD1P3AX array_255___i329 (.D(array_0__7__N_3769[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[214] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i329.GSR = "ENABLED";
    FD1P3AX array_255___i330 (.D(array_0__7__N_3769[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[214] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i330.GSR = "ENABLED";
    FD1P3AX array_255___i331 (.D(array_0__7__N_3769[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[214] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i331.GSR = "ENABLED";
    FD1P3AX array_255___i332 (.D(array_0__7__N_3769[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[214] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i332.GSR = "ENABLED";
    FD1P3AX array_255___i333 (.D(array_0__7__N_3769[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[214] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i333.GSR = "ENABLED";
    FD1P3AX array_255___i334 (.D(array_0__7__N_3769[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[214] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i334.GSR = "ENABLED";
    FD1P3AX array_255___i335 (.D(array_0__7__N_3769[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[214] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i335.GSR = "ENABLED";
    FD1P3AX array_255___i336 (.D(array_0__7__N_3769[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[214] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i336.GSR = "ENABLED";
    FD1P3AX array_255___i337 (.D(array_0__7__N_3761[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[213] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i337.GSR = "ENABLED";
    FD1P3AX array_255___i338 (.D(array_0__7__N_3761[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[213] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i338.GSR = "ENABLED";
    FD1P3AX array_255___i339 (.D(array_0__7__N_3761[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[213] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i339.GSR = "ENABLED";
    FD1P3AX array_255___i340 (.D(array_0__7__N_3761[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[213] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i340.GSR = "ENABLED";
    FD1P3AX array_255___i341 (.D(array_0__7__N_3761[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[213] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i341.GSR = "ENABLED";
    FD1P3AX array_255___i342 (.D(array_0__7__N_3761[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[213] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i342.GSR = "ENABLED";
    FD1P3AX array_255___i343 (.D(array_0__7__N_3761[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[213] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i343.GSR = "ENABLED";
    FD1P3AX array_255___i344 (.D(array_0__7__N_3761[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[213] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i344.GSR = "ENABLED";
    FD1P3AX array_255___i345 (.D(array_0__7__N_3753[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[212] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i345.GSR = "ENABLED";
    FD1P3AX array_255___i346 (.D(array_0__7__N_3753[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[212] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i346.GSR = "ENABLED";
    FD1P3AX array_255___i347 (.D(array_0__7__N_3753[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[212] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i347.GSR = "ENABLED";
    FD1P3AX array_255___i348 (.D(array_0__7__N_3753[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[212] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i348.GSR = "ENABLED";
    FD1P3AX array_255___i349 (.D(array_0__7__N_3753[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[212] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i349.GSR = "ENABLED";
    FD1P3AX array_255___i350 (.D(array_0__7__N_3753[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[212] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i350.GSR = "ENABLED";
    FD1P3AX array_255___i351 (.D(array_0__7__N_3753[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[212] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i351.GSR = "ENABLED";
    FD1P3AX array_255___i352 (.D(array_0__7__N_3753[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[212] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i352.GSR = "ENABLED";
    FD1P3AX array_255___i353 (.D(array_0__7__N_3745[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[211] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i353.GSR = "ENABLED";
    FD1P3AX array_255___i354 (.D(array_0__7__N_3745[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[211] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i354.GSR = "ENABLED";
    FD1P3AX array_255___i355 (.D(array_0__7__N_3745[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[211] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i355.GSR = "ENABLED";
    FD1P3AX array_255___i356 (.D(array_0__7__N_3745[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[211] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i356.GSR = "ENABLED";
    FD1P3AX array_255___i357 (.D(array_0__7__N_3745[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[211] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i357.GSR = "ENABLED";
    FD1P3AX array_255___i358 (.D(array_0__7__N_3745[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[211] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i358.GSR = "ENABLED";
    FD1P3AX array_255___i359 (.D(array_0__7__N_3745[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[211] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i359.GSR = "ENABLED";
    FD1P3AX array_255___i360 (.D(array_0__7__N_3745[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[211] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i360.GSR = "ENABLED";
    FD1P3AX array_255___i361 (.D(array_0__7__N_3737[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[210] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i361.GSR = "ENABLED";
    FD1P3AX array_255___i362 (.D(array_0__7__N_3737[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[210] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i362.GSR = "ENABLED";
    FD1P3AX array_255___i363 (.D(array_0__7__N_3737[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[210] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i363.GSR = "ENABLED";
    FD1P3AX array_255___i364 (.D(array_0__7__N_3737[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[210] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i364.GSR = "ENABLED";
    FD1P3AX array_255___i365 (.D(array_0__7__N_3737[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[210] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i365.GSR = "ENABLED";
    FD1P3AX array_255___i366 (.D(array_0__7__N_3737[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[210] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i366.GSR = "ENABLED";
    FD1P3AX array_255___i367 (.D(array_0__7__N_3737[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[210] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i367.GSR = "ENABLED";
    FD1P3AX array_255___i368 (.D(array_0__7__N_3737[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[210] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i368.GSR = "ENABLED";
    FD1P3AX array_255___i369 (.D(array_0__7__N_3729[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[209] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i369.GSR = "ENABLED";
    FD1P3AX array_255___i370 (.D(array_0__7__N_3729[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[209] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i370.GSR = "ENABLED";
    FD1P3AX array_255___i371 (.D(array_0__7__N_3729[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[209] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i371.GSR = "ENABLED";
    FD1P3AX array_255___i372 (.D(array_0__7__N_3729[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[209] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i372.GSR = "ENABLED";
    FD1P3AX array_255___i373 (.D(array_0__7__N_3729[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[209] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i373.GSR = "ENABLED";
    FD1P3AX array_255___i374 (.D(array_0__7__N_3729[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[209] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i374.GSR = "ENABLED";
    FD1P3AX array_255___i375 (.D(array_0__7__N_3729[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[209] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i375.GSR = "ENABLED";
    FD1P3AX array_255___i376 (.D(array_0__7__N_3729[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[209] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i376.GSR = "ENABLED";
    FD1P3AX array_255___i377 (.D(array_0__7__N_3721[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[208] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i377.GSR = "ENABLED";
    FD1P3AX array_255___i378 (.D(array_0__7__N_3721[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[208] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i378.GSR = "ENABLED";
    FD1P3AX array_255___i379 (.D(array_0__7__N_3721[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[208] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i379.GSR = "ENABLED";
    FD1P3AX array_255___i380 (.D(array_0__7__N_3721[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[208] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i380.GSR = "ENABLED";
    FD1P3AX array_255___i381 (.D(array_0__7__N_3721[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[208] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i381.GSR = "ENABLED";
    FD1P3AX array_255___i382 (.D(array_0__7__N_3721[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[208] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i382.GSR = "ENABLED";
    FD1P3AX array_255___i383 (.D(array_0__7__N_3721[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[208] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i383.GSR = "ENABLED";
    FD1P3AX array_255___i384 (.D(array_0__7__N_3721[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[208] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i384.GSR = "ENABLED";
    FD1P3AX array_255___i385 (.D(array_0__7__N_3713[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[207] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i385.GSR = "ENABLED";
    FD1P3AX array_255___i386 (.D(array_0__7__N_3713[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[207] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i386.GSR = "ENABLED";
    FD1P3AX array_255___i387 (.D(array_0__7__N_3713[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[207] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i387.GSR = "ENABLED";
    FD1P3AX array_255___i388 (.D(array_0__7__N_3713[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[207] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i388.GSR = "ENABLED";
    FD1P3AX array_255___i389 (.D(array_0__7__N_3713[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[207] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i389.GSR = "ENABLED";
    FD1P3AX array_255___i390 (.D(array_0__7__N_3713[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[207] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i390.GSR = "ENABLED";
    FD1P3AX array_255___i391 (.D(array_0__7__N_3713[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[207] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i391.GSR = "ENABLED";
    FD1P3AX array_255___i392 (.D(array_0__7__N_3713[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[207] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i392.GSR = "ENABLED";
    FD1P3AX array_255___i393 (.D(array_0__7__N_3705[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[206] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i393.GSR = "ENABLED";
    FD1P3AX array_255___i394 (.D(array_0__7__N_3705[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[206] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i394.GSR = "ENABLED";
    FD1P3AX array_255___i395 (.D(array_0__7__N_3705[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[206] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i395.GSR = "ENABLED";
    FD1P3AX array_255___i396 (.D(array_0__7__N_3705[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[206] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i396.GSR = "ENABLED";
    FD1P3AX array_255___i397 (.D(array_0__7__N_3705[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[206] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i397.GSR = "ENABLED";
    FD1P3AX array_255___i398 (.D(array_0__7__N_3705[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[206] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i398.GSR = "ENABLED";
    FD1P3AX array_255___i399 (.D(array_0__7__N_3705[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[206] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i399.GSR = "ENABLED";
    FD1P3AX array_255___i400 (.D(array_0__7__N_3705[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[206] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i400.GSR = "ENABLED";
    FD1P3AX array_255___i401 (.D(array_0__7__N_3697[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[205] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i401.GSR = "ENABLED";
    FD1P3AX array_255___i402 (.D(array_0__7__N_3697[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[205] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i402.GSR = "ENABLED";
    FD1P3AX array_255___i403 (.D(array_0__7__N_3697[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[205] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i403.GSR = "ENABLED";
    FD1P3AX array_255___i404 (.D(array_0__7__N_3697[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[205] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i404.GSR = "ENABLED";
    FD1P3AX array_255___i405 (.D(array_0__7__N_3697[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[205] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i405.GSR = "ENABLED";
    FD1P3AX array_255___i406 (.D(array_0__7__N_3697[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[205] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i406.GSR = "ENABLED";
    FD1P3AX array_255___i407 (.D(array_0__7__N_3697[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[205] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i407.GSR = "ENABLED";
    FD1P3AX array_255___i408 (.D(array_0__7__N_3697[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[205] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i408.GSR = "ENABLED";
    FD1P3AX array_255___i409 (.D(array_0__7__N_3689[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[204] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i409.GSR = "ENABLED";
    FD1P3AX array_255___i410 (.D(array_0__7__N_3689[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[204] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i410.GSR = "ENABLED";
    FD1P3AX array_255___i411 (.D(array_0__7__N_3689[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[204] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i411.GSR = "ENABLED";
    FD1P3AX array_255___i412 (.D(array_0__7__N_3689[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[204] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i412.GSR = "ENABLED";
    FD1P3AX array_255___i413 (.D(array_0__7__N_3689[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[204] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i413.GSR = "ENABLED";
    FD1P3AX array_255___i414 (.D(array_0__7__N_3689[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[204] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i414.GSR = "ENABLED";
    FD1P3AX array_255___i415 (.D(array_0__7__N_3689[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[204] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i415.GSR = "ENABLED";
    FD1P3AX array_255___i416 (.D(array_0__7__N_3689[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[204] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i416.GSR = "ENABLED";
    FD1P3AX array_255___i417 (.D(array_0__7__N_3681[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[203] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i417.GSR = "ENABLED";
    FD1P3AX array_255___i418 (.D(array_0__7__N_3681[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[203] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i418.GSR = "ENABLED";
    FD1P3AX array_255___i419 (.D(array_0__7__N_3681[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[203] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i419.GSR = "ENABLED";
    FD1P3AX array_255___i420 (.D(array_0__7__N_3681[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[203] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i420.GSR = "ENABLED";
    FD1P3AX array_255___i421 (.D(array_0__7__N_3681[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[203] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i421.GSR = "ENABLED";
    FD1P3AX array_255___i422 (.D(array_0__7__N_3681[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[203] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i422.GSR = "ENABLED";
    FD1P3AX array_255___i423 (.D(array_0__7__N_3681[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[203] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i423.GSR = "ENABLED";
    FD1P3AX array_255___i424 (.D(array_0__7__N_3681[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[203] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i424.GSR = "ENABLED";
    FD1P3AX array_255___i425 (.D(array_0__7__N_3673[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[202] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i425.GSR = "ENABLED";
    FD1P3AX array_255___i426 (.D(array_0__7__N_3673[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[202] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i426.GSR = "ENABLED";
    FD1P3AX array_255___i427 (.D(array_0__7__N_3673[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[202] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i427.GSR = "ENABLED";
    FD1P3AX array_255___i428 (.D(array_0__7__N_3673[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[202] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i428.GSR = "ENABLED";
    FD1P3AX array_255___i429 (.D(array_0__7__N_3673[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[202] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i429.GSR = "ENABLED";
    FD1P3AX array_255___i430 (.D(array_0__7__N_3673[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[202] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i430.GSR = "ENABLED";
    FD1P3AX array_255___i431 (.D(array_0__7__N_3673[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[202] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i431.GSR = "ENABLED";
    FD1P3AX array_255___i432 (.D(array_0__7__N_3673[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[202] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i432.GSR = "ENABLED";
    FD1P3AX array_255___i433 (.D(array_0__7__N_3665[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[201] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i433.GSR = "ENABLED";
    FD1P3AX array_255___i434 (.D(array_0__7__N_3665[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[201] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i434.GSR = "ENABLED";
    FD1P3AX array_255___i435 (.D(array_0__7__N_3665[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[201] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i435.GSR = "ENABLED";
    FD1P3AX array_255___i436 (.D(array_0__7__N_3665[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[201] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i436.GSR = "ENABLED";
    FD1P3AX array_255___i437 (.D(array_0__7__N_3665[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[201] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i437.GSR = "ENABLED";
    FD1P3AX array_255___i438 (.D(array_0__7__N_3665[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[201] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i438.GSR = "ENABLED";
    FD1P3AX array_255___i439 (.D(array_0__7__N_3665[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[201] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i439.GSR = "ENABLED";
    FD1P3AX array_255___i440 (.D(array_0__7__N_3665[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[201] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i440.GSR = "ENABLED";
    FD1P3AX array_255___i441 (.D(array_0__7__N_3657[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[200] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i441.GSR = "ENABLED";
    FD1P3AX array_255___i442 (.D(array_0__7__N_3657[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[200] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i442.GSR = "ENABLED";
    FD1P3AX array_255___i443 (.D(array_0__7__N_3657[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[200] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i443.GSR = "ENABLED";
    FD1P3AX array_255___i444 (.D(array_0__7__N_3657[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[200] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i444.GSR = "ENABLED";
    FD1P3AX array_255___i445 (.D(array_0__7__N_3657[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[200] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i445.GSR = "ENABLED";
    FD1P3AX array_255___i446 (.D(array_0__7__N_3657[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[200] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i446.GSR = "ENABLED";
    FD1P3AX array_255___i447 (.D(array_0__7__N_3657[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[200] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i447.GSR = "ENABLED";
    FD1P3AX array_255___i448 (.D(array_0__7__N_3657[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[200] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i448.GSR = "ENABLED";
    FD1P3AX array_255___i449 (.D(array_0__7__N_3649[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[199] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i449.GSR = "ENABLED";
    FD1P3AX array_255___i450 (.D(array_0__7__N_3649[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[199] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i450.GSR = "ENABLED";
    FD1P3AX array_255___i451 (.D(array_0__7__N_3649[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[199] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i451.GSR = "ENABLED";
    FD1P3AX array_255___i452 (.D(array_0__7__N_3649[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[199] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i452.GSR = "ENABLED";
    FD1P3AX array_255___i453 (.D(array_0__7__N_3649[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[199] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i453.GSR = "ENABLED";
    FD1P3AX array_255___i454 (.D(array_0__7__N_3649[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[199] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i454.GSR = "ENABLED";
    FD1P3AX array_255___i455 (.D(array_0__7__N_3649[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[199] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i455.GSR = "ENABLED";
    FD1P3AX array_255___i456 (.D(array_0__7__N_3649[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[199] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i456.GSR = "ENABLED";
    FD1P3AX array_255___i457 (.D(array_0__7__N_3641[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[198] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i457.GSR = "ENABLED";
    FD1P3AX array_255___i458 (.D(array_0__7__N_3641[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[198] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i458.GSR = "ENABLED";
    FD1P3AX array_255___i459 (.D(array_0__7__N_3641[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[198] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i459.GSR = "ENABLED";
    FD1P3AX array_255___i460 (.D(array_0__7__N_3641[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[198] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i460.GSR = "ENABLED";
    FD1P3AX array_255___i461 (.D(array_0__7__N_3641[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[198] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i461.GSR = "ENABLED";
    FD1P3AX array_255___i462 (.D(array_0__7__N_3641[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[198] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i462.GSR = "ENABLED";
    FD1P3AX array_255___i463 (.D(array_0__7__N_3641[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[198] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i463.GSR = "ENABLED";
    FD1P3AX array_255___i464 (.D(array_0__7__N_3641[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[198] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i464.GSR = "ENABLED";
    FD1P3AX array_255___i465 (.D(array_0__7__N_3633[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[197] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i465.GSR = "ENABLED";
    FD1P3AX array_255___i466 (.D(array_0__7__N_3633[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[197] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i466.GSR = "ENABLED";
    FD1P3AX array_255___i467 (.D(array_0__7__N_3633[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[197] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i467.GSR = "ENABLED";
    FD1P3AX array_255___i468 (.D(array_0__7__N_3633[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[197] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i468.GSR = "ENABLED";
    FD1P3AX array_255___i469 (.D(array_0__7__N_3633[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[197] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i469.GSR = "ENABLED";
    FD1P3AX array_255___i470 (.D(array_0__7__N_3633[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[197] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i470.GSR = "ENABLED";
    FD1P3AX array_255___i471 (.D(array_0__7__N_3633[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[197] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i471.GSR = "ENABLED";
    FD1P3AX array_255___i472 (.D(array_0__7__N_3633[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[197] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i472.GSR = "ENABLED";
    FD1P3AX array_255___i473 (.D(array_0__7__N_3625[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[196] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i473.GSR = "ENABLED";
    FD1P3AX array_255___i474 (.D(array_0__7__N_3625[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[196] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i474.GSR = "ENABLED";
    FD1P3AX array_255___i475 (.D(array_0__7__N_3625[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[196] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i475.GSR = "ENABLED";
    FD1P3AX array_255___i476 (.D(array_0__7__N_3625[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[196] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i476.GSR = "ENABLED";
    FD1P3AX array_255___i477 (.D(array_0__7__N_3625[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[196] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i477.GSR = "ENABLED";
    FD1P3AX array_255___i478 (.D(array_0__7__N_3625[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[196] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i478.GSR = "ENABLED";
    FD1P3AX array_255___i479 (.D(array_0__7__N_3625[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[196] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i479.GSR = "ENABLED";
    FD1P3AX array_255___i480 (.D(array_0__7__N_3625[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[196] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i480.GSR = "ENABLED";
    FD1P3AX array_255___i481 (.D(array_0__7__N_3617[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[195] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i481.GSR = "ENABLED";
    FD1P3AX array_255___i482 (.D(array_0__7__N_3617[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[195] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i482.GSR = "ENABLED";
    FD1P3AX array_255___i483 (.D(array_0__7__N_3617[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[195] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i483.GSR = "ENABLED";
    FD1P3AX array_255___i484 (.D(array_0__7__N_3617[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[195] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i484.GSR = "ENABLED";
    FD1P3AX array_255___i485 (.D(array_0__7__N_3617[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[195] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i485.GSR = "ENABLED";
    FD1P3AX array_255___i486 (.D(array_0__7__N_3617[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[195] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i486.GSR = "ENABLED";
    FD1P3AX array_255___i487 (.D(array_0__7__N_3617[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[195] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i487.GSR = "ENABLED";
    FD1P3AX array_255___i488 (.D(array_0__7__N_3617[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[195] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i488.GSR = "ENABLED";
    FD1P3AX array_255___i489 (.D(array_0__7__N_3609[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[194] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i489.GSR = "ENABLED";
    FD1P3AX array_255___i490 (.D(array_0__7__N_3609[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[194] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i490.GSR = "ENABLED";
    FD1P3AX array_255___i491 (.D(array_0__7__N_3609[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[194] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i491.GSR = "ENABLED";
    FD1P3AX array_255___i492 (.D(array_0__7__N_3609[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[194] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i492.GSR = "ENABLED";
    FD1P3AX array_255___i493 (.D(array_0__7__N_3609[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[194] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i493.GSR = "ENABLED";
    FD1P3AX array_255___i494 (.D(array_0__7__N_3609[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[194] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i494.GSR = "ENABLED";
    FD1P3AX array_255___i495 (.D(array_0__7__N_3609[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[194] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i495.GSR = "ENABLED";
    FD1P3AX array_255___i496 (.D(array_0__7__N_3609[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[194] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i496.GSR = "ENABLED";
    FD1P3AX array_255___i497 (.D(array_0__7__N_3601[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[193] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i497.GSR = "ENABLED";
    FD1P3AX array_255___i498 (.D(array_0__7__N_3601[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[193] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i498.GSR = "ENABLED";
    FD1P3AX array_255___i499 (.D(array_0__7__N_3601[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[193] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i499.GSR = "ENABLED";
    FD1P3AX array_255___i500 (.D(array_0__7__N_3601[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[193] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i500.GSR = "ENABLED";
    FD1P3AX array_255___i501 (.D(array_0__7__N_3601[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[193] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i501.GSR = "ENABLED";
    FD1P3AX array_255___i502 (.D(array_0__7__N_3601[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[193] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i502.GSR = "ENABLED";
    FD1P3AX array_255___i503 (.D(array_0__7__N_3601[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[193] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i503.GSR = "ENABLED";
    FD1P3AX array_255___i504 (.D(array_0__7__N_3601[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[193] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i504.GSR = "ENABLED";
    FD1P3AX array_255___i505 (.D(array_0__7__N_3593[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[192] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i505.GSR = "ENABLED";
    FD1P3AX array_255___i506 (.D(array_0__7__N_3593[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[192] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i506.GSR = "ENABLED";
    FD1P3AX array_255___i507 (.D(array_0__7__N_3593[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[192] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i507.GSR = "ENABLED";
    FD1P3AX array_255___i508 (.D(array_0__7__N_3593[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[192] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i508.GSR = "ENABLED";
    FD1P3AX array_255___i509 (.D(array_0__7__N_3593[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[192] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i509.GSR = "ENABLED";
    FD1P3AX array_255___i510 (.D(array_0__7__N_3593[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[192] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i510.GSR = "ENABLED";
    FD1P3AX array_255___i511 (.D(array_0__7__N_3593[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[192] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i511.GSR = "ENABLED";
    FD1P3AX array_255___i512 (.D(array_0__7__N_3593[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[192] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i512.GSR = "ENABLED";
    FD1P3AX array_255___i513 (.D(array_0__7__N_3585[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[191] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i513.GSR = "ENABLED";
    FD1P3AX array_255___i514 (.D(array_0__7__N_3585[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[191] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i514.GSR = "ENABLED";
    FD1P3AX array_255___i515 (.D(array_0__7__N_3585[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[191] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i515.GSR = "ENABLED";
    FD1P3AX array_255___i516 (.D(array_0__7__N_3585[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[191] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i516.GSR = "ENABLED";
    FD1P3AX array_255___i517 (.D(array_0__7__N_3585[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[191] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i517.GSR = "ENABLED";
    FD1P3AX array_255___i518 (.D(array_0__7__N_3585[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[191] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i518.GSR = "ENABLED";
    FD1P3AX array_255___i519 (.D(array_0__7__N_3585[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[191] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i519.GSR = "ENABLED";
    FD1P3AX array_255___i520 (.D(array_0__7__N_3585[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[191] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i520.GSR = "ENABLED";
    FD1P3AX array_255___i521 (.D(array_0__7__N_3577[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[190] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i521.GSR = "ENABLED";
    FD1P3AX array_255___i522 (.D(array_0__7__N_3577[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[190] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i522.GSR = "ENABLED";
    FD1P3AX array_255___i523 (.D(array_0__7__N_3577[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[190] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i523.GSR = "ENABLED";
    FD1P3AX array_255___i524 (.D(array_0__7__N_3577[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[190] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i524.GSR = "ENABLED";
    FD1P3AX array_255___i525 (.D(array_0__7__N_3577[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[190] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i525.GSR = "ENABLED";
    FD1P3AX array_255___i526 (.D(array_0__7__N_3577[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[190] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i526.GSR = "ENABLED";
    FD1P3AX array_255___i527 (.D(array_0__7__N_3577[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[190] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i527.GSR = "ENABLED";
    FD1P3AX array_255___i528 (.D(array_0__7__N_3577[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[190] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i528.GSR = "ENABLED";
    FD1P3AX array_255___i529 (.D(array_0__7__N_3569[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[189] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i529.GSR = "ENABLED";
    FD1P3AX array_255___i530 (.D(array_0__7__N_3569[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[189] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i530.GSR = "ENABLED";
    FD1P3AX array_255___i531 (.D(array_0__7__N_3569[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[189] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i531.GSR = "ENABLED";
    FD1P3AX array_255___i532 (.D(array_0__7__N_3569[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[189] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i532.GSR = "ENABLED";
    FD1P3AX array_255___i533 (.D(array_0__7__N_3569[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[189] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i533.GSR = "ENABLED";
    FD1P3AX array_255___i534 (.D(array_0__7__N_3569[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[189] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i534.GSR = "ENABLED";
    FD1P3AX array_255___i535 (.D(array_0__7__N_3569[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[189] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i535.GSR = "ENABLED";
    FD1P3AX array_255___i536 (.D(array_0__7__N_3569[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[189] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i536.GSR = "ENABLED";
    FD1P3AX array_255___i537 (.D(array_0__7__N_3561[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[188] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i537.GSR = "ENABLED";
    FD1P3AX array_255___i538 (.D(array_0__7__N_3561[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[188] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i538.GSR = "ENABLED";
    FD1P3AX array_255___i539 (.D(array_0__7__N_3561[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[188] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i539.GSR = "ENABLED";
    FD1P3AX array_255___i540 (.D(array_0__7__N_3561[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[188] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i540.GSR = "ENABLED";
    FD1P3AX array_255___i541 (.D(array_0__7__N_3561[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[188] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i541.GSR = "ENABLED";
    FD1P3AX array_255___i542 (.D(array_0__7__N_3561[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[188] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i542.GSR = "ENABLED";
    FD1P3AX array_255___i543 (.D(array_0__7__N_3561[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[188] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i543.GSR = "ENABLED";
    FD1P3AX array_255___i544 (.D(array_0__7__N_3561[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[188] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i544.GSR = "ENABLED";
    FD1P3AX array_255___i545 (.D(array_0__7__N_3553[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[187] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i545.GSR = "ENABLED";
    FD1P3AX array_255___i546 (.D(array_0__7__N_3553[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[187] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i546.GSR = "ENABLED";
    FD1P3AX array_255___i547 (.D(array_0__7__N_3553[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[187] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i547.GSR = "ENABLED";
    FD1P3AX array_255___i548 (.D(array_0__7__N_3553[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[187] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i548.GSR = "ENABLED";
    FD1P3AX array_255___i549 (.D(array_0__7__N_3553[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[187] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i549.GSR = "ENABLED";
    FD1P3AX array_255___i550 (.D(array_0__7__N_3553[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[187] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i550.GSR = "ENABLED";
    FD1P3AX array_255___i551 (.D(array_0__7__N_3553[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[187] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i551.GSR = "ENABLED";
    FD1P3AX array_255___i552 (.D(array_0__7__N_3553[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[187] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i552.GSR = "ENABLED";
    FD1P3AX array_255___i553 (.D(array_0__7__N_3545[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[186] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i553.GSR = "ENABLED";
    FD1P3AX array_255___i554 (.D(array_0__7__N_3545[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[186] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i554.GSR = "ENABLED";
    FD1P3AX array_255___i555 (.D(array_0__7__N_3545[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[186] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i555.GSR = "ENABLED";
    FD1P3AX array_255___i556 (.D(array_0__7__N_3545[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[186] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i556.GSR = "ENABLED";
    FD1P3AX array_255___i557 (.D(array_0__7__N_3545[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[186] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i557.GSR = "ENABLED";
    FD1P3AX array_255___i558 (.D(array_0__7__N_3545[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[186] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i558.GSR = "ENABLED";
    FD1P3AX array_255___i559 (.D(array_0__7__N_3545[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[186] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i559.GSR = "ENABLED";
    FD1P3AX array_255___i560 (.D(array_0__7__N_3545[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[186] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i560.GSR = "ENABLED";
    FD1P3AX array_255___i561 (.D(array_0__7__N_3537[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[185] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i561.GSR = "ENABLED";
    FD1P3AX array_255___i562 (.D(array_0__7__N_3537[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[185] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i562.GSR = "ENABLED";
    FD1P3AX array_255___i563 (.D(array_0__7__N_3537[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[185] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i563.GSR = "ENABLED";
    FD1P3AX array_255___i564 (.D(array_0__7__N_3537[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[185] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i564.GSR = "ENABLED";
    FD1P3AX array_255___i565 (.D(array_0__7__N_3537[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[185] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i565.GSR = "ENABLED";
    FD1P3AX array_255___i566 (.D(array_0__7__N_3537[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[185] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i566.GSR = "ENABLED";
    FD1P3AX array_255___i567 (.D(array_0__7__N_3537[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[185] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i567.GSR = "ENABLED";
    FD1P3AX array_255___i568 (.D(array_0__7__N_3537[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[185] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i568.GSR = "ENABLED";
    FD1P3AX array_255___i569 (.D(array_0__7__N_3529[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[184] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i569.GSR = "ENABLED";
    FD1P3AX array_255___i570 (.D(array_0__7__N_3529[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[184] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i570.GSR = "ENABLED";
    FD1P3AX array_255___i571 (.D(array_0__7__N_3529[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[184] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i571.GSR = "ENABLED";
    FD1P3AX array_255___i572 (.D(array_0__7__N_3529[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[184] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i572.GSR = "ENABLED";
    FD1P3AX array_255___i573 (.D(array_0__7__N_3529[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[184] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i573.GSR = "ENABLED";
    FD1P3AX array_255___i574 (.D(array_0__7__N_3529[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[184] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i574.GSR = "ENABLED";
    FD1P3AX array_255___i575 (.D(array_0__7__N_3529[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[184] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i575.GSR = "ENABLED";
    FD1P3AX array_255___i576 (.D(array_0__7__N_3529[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[184] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i576.GSR = "ENABLED";
    FD1P3AX array_255___i577 (.D(array_0__7__N_3521[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[183] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i577.GSR = "ENABLED";
    FD1P3AX array_255___i578 (.D(array_0__7__N_3521[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[183] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i578.GSR = "ENABLED";
    FD1P3AX array_255___i579 (.D(array_0__7__N_3521[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[183] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i579.GSR = "ENABLED";
    FD1P3AX array_255___i580 (.D(array_0__7__N_3521[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[183] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i580.GSR = "ENABLED";
    FD1P3AX array_255___i581 (.D(array_0__7__N_3521[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[183] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i581.GSR = "ENABLED";
    FD1P3AX array_255___i582 (.D(array_0__7__N_3521[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[183] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i582.GSR = "ENABLED";
    FD1P3AX array_255___i583 (.D(array_0__7__N_3521[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[183] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i583.GSR = "ENABLED";
    FD1P3AX array_255___i584 (.D(array_0__7__N_3521[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[183] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i584.GSR = "ENABLED";
    FD1P3AX array_255___i585 (.D(array_0__7__N_3513[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[182] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i585.GSR = "ENABLED";
    FD1P3AX array_255___i586 (.D(array_0__7__N_3513[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[182] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i586.GSR = "ENABLED";
    FD1P3AX array_255___i587 (.D(array_0__7__N_3513[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[182] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i587.GSR = "ENABLED";
    FD1P3AX array_255___i588 (.D(array_0__7__N_3513[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[182] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i588.GSR = "ENABLED";
    FD1P3AX array_255___i589 (.D(array_0__7__N_3513[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[182] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i589.GSR = "ENABLED";
    FD1P3AX array_255___i590 (.D(array_0__7__N_3513[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[182] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i590.GSR = "ENABLED";
    FD1P3AX array_255___i591 (.D(array_0__7__N_3513[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[182] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i591.GSR = "ENABLED";
    FD1P3AX array_255___i592 (.D(array_0__7__N_3513[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[182] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i592.GSR = "ENABLED";
    FD1P3AX array_255___i593 (.D(array_0__7__N_3505[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[181] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i593.GSR = "ENABLED";
    FD1P3AX array_255___i594 (.D(array_0__7__N_3505[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[181] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i594.GSR = "ENABLED";
    FD1P3AX array_255___i595 (.D(array_0__7__N_3505[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[181] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i595.GSR = "ENABLED";
    FD1P3AX array_255___i596 (.D(array_0__7__N_3505[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[181] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i596.GSR = "ENABLED";
    FD1P3AX array_255___i597 (.D(array_0__7__N_3505[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[181] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i597.GSR = "ENABLED";
    FD1P3AX array_255___i598 (.D(array_0__7__N_3505[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[181] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i598.GSR = "ENABLED";
    FD1P3AX array_255___i599 (.D(array_0__7__N_3505[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[181] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i599.GSR = "ENABLED";
    FD1P3AX array_255___i600 (.D(array_0__7__N_3505[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[181] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i600.GSR = "ENABLED";
    FD1P3AX array_255___i601 (.D(array_0__7__N_3497[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[180] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i601.GSR = "ENABLED";
    FD1P3AX array_255___i602 (.D(array_0__7__N_3497[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[180] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i602.GSR = "ENABLED";
    FD1P3AX array_255___i603 (.D(array_0__7__N_3497[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[180] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i603.GSR = "ENABLED";
    FD1P3AX array_255___i604 (.D(array_0__7__N_3497[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[180] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i604.GSR = "ENABLED";
    FD1P3AX array_255___i605 (.D(array_0__7__N_3497[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[180] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i605.GSR = "ENABLED";
    FD1P3AX array_255___i606 (.D(array_0__7__N_3497[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[180] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i606.GSR = "ENABLED";
    FD1P3AX array_255___i607 (.D(array_0__7__N_3497[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[180] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i607.GSR = "ENABLED";
    FD1P3AX array_255___i608 (.D(array_0__7__N_3497[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[180] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i608.GSR = "ENABLED";
    FD1P3AX array_255___i609 (.D(array_0__7__N_3489[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[179] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i609.GSR = "ENABLED";
    FD1P3AX array_255___i610 (.D(array_0__7__N_3489[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[179] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i610.GSR = "ENABLED";
    FD1P3AX array_255___i611 (.D(array_0__7__N_3489[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[179] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i611.GSR = "ENABLED";
    FD1P3AX array_255___i612 (.D(array_0__7__N_3489[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[179] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i612.GSR = "ENABLED";
    FD1P3AX array_255___i613 (.D(array_0__7__N_3489[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[179] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i613.GSR = "ENABLED";
    FD1P3AX array_255___i614 (.D(array_0__7__N_3489[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[179] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i614.GSR = "ENABLED";
    FD1P3AX array_255___i615 (.D(array_0__7__N_3489[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[179] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i615.GSR = "ENABLED";
    FD1P3AX array_255___i616 (.D(array_0__7__N_3489[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[179] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i616.GSR = "ENABLED";
    FD1P3AX array_255___i617 (.D(array_0__7__N_3481[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[178] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i617.GSR = "ENABLED";
    FD1P3AX array_255___i618 (.D(array_0__7__N_3481[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[178] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i618.GSR = "ENABLED";
    FD1P3AX array_255___i619 (.D(array_0__7__N_3481[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[178] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i619.GSR = "ENABLED";
    FD1P3AX array_255___i620 (.D(array_0__7__N_3481[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[178] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i620.GSR = "ENABLED";
    FD1P3AX array_255___i621 (.D(array_0__7__N_3481[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[178] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i621.GSR = "ENABLED";
    FD1P3AX array_255___i622 (.D(array_0__7__N_3481[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[178] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i622.GSR = "ENABLED";
    FD1P3AX array_255___i623 (.D(array_0__7__N_3481[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[178] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i623.GSR = "ENABLED";
    FD1P3AX array_255___i624 (.D(array_0__7__N_3481[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[178] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i624.GSR = "ENABLED";
    FD1P3AX array_255___i625 (.D(array_0__7__N_3473[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[177] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i625.GSR = "ENABLED";
    FD1P3AX array_255___i626 (.D(array_0__7__N_3473[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[177] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i626.GSR = "ENABLED";
    FD1P3AX array_255___i627 (.D(array_0__7__N_3473[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[177] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i627.GSR = "ENABLED";
    FD1P3AX array_255___i628 (.D(array_0__7__N_3473[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[177] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i628.GSR = "ENABLED";
    FD1P3AX array_255___i629 (.D(array_0__7__N_3473[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[177] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i629.GSR = "ENABLED";
    FD1P3AX array_255___i630 (.D(array_0__7__N_3473[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[177] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i630.GSR = "ENABLED";
    FD1P3AX array_255___i631 (.D(array_0__7__N_3473[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[177] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i631.GSR = "ENABLED";
    FD1P3AX array_255___i632 (.D(array_0__7__N_3473[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[177] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i632.GSR = "ENABLED";
    FD1P3AX array_255___i633 (.D(array_0__7__N_3465[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[176] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i633.GSR = "ENABLED";
    FD1P3AX array_255___i634 (.D(array_0__7__N_3465[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[176] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i634.GSR = "ENABLED";
    FD1P3AX array_255___i635 (.D(array_0__7__N_3465[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[176] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i635.GSR = "ENABLED";
    FD1P3AX array_255___i636 (.D(array_0__7__N_3465[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[176] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i636.GSR = "ENABLED";
    FD1P3AX array_255___i637 (.D(array_0__7__N_3465[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[176] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i637.GSR = "ENABLED";
    FD1P3AX array_255___i638 (.D(array_0__7__N_3465[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[176] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i638.GSR = "ENABLED";
    FD1P3AX array_255___i639 (.D(array_0__7__N_3465[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[176] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i639.GSR = "ENABLED";
    FD1P3AX array_255___i640 (.D(array_0__7__N_3465[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[176] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i640.GSR = "ENABLED";
    FD1P3AX array_255___i641 (.D(array_0__7__N_3457[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[175] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i641.GSR = "ENABLED";
    FD1P3AX array_255___i642 (.D(array_0__7__N_3457[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[175] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i642.GSR = "ENABLED";
    FD1P3AX array_255___i643 (.D(array_0__7__N_3457[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[175] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i643.GSR = "ENABLED";
    FD1P3AX array_255___i644 (.D(array_0__7__N_3457[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[175] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i644.GSR = "ENABLED";
    FD1P3AX array_255___i645 (.D(array_0__7__N_3457[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[175] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i645.GSR = "ENABLED";
    FD1P3AX array_255___i646 (.D(array_0__7__N_3457[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[175] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i646.GSR = "ENABLED";
    FD1P3AX array_255___i647 (.D(array_0__7__N_3457[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[175] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i647.GSR = "ENABLED";
    FD1P3AX array_255___i648 (.D(array_0__7__N_3457[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[175] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i648.GSR = "ENABLED";
    FD1P3AX array_255___i649 (.D(array_0__7__N_3449[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[174] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i649.GSR = "ENABLED";
    FD1P3AX array_255___i650 (.D(array_0__7__N_3449[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[174] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i650.GSR = "ENABLED";
    FD1P3AX array_255___i651 (.D(array_0__7__N_3449[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[174] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i651.GSR = "ENABLED";
    FD1P3AX array_255___i652 (.D(array_0__7__N_3449[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[174] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i652.GSR = "ENABLED";
    FD1P3AX array_255___i653 (.D(array_0__7__N_3449[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[174] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i653.GSR = "ENABLED";
    FD1P3AX array_255___i654 (.D(array_0__7__N_3449[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[174] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i654.GSR = "ENABLED";
    FD1P3AX array_255___i655 (.D(array_0__7__N_3449[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[174] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i655.GSR = "ENABLED";
    FD1P3AX array_255___i656 (.D(array_0__7__N_3449[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[174] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i656.GSR = "ENABLED";
    FD1P3AX array_255___i657 (.D(array_0__7__N_3441[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[173] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i657.GSR = "ENABLED";
    FD1P3AX array_255___i658 (.D(array_0__7__N_3441[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[173] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i658.GSR = "ENABLED";
    FD1P3AX array_255___i659 (.D(array_0__7__N_3441[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[173] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i659.GSR = "ENABLED";
    FD1P3AX array_255___i660 (.D(array_0__7__N_3441[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[173] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i660.GSR = "ENABLED";
    FD1P3AX array_255___i661 (.D(array_0__7__N_3441[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[173] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i661.GSR = "ENABLED";
    FD1P3AX array_255___i662 (.D(array_0__7__N_3441[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[173] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i662.GSR = "ENABLED";
    FD1P3AX array_255___i663 (.D(array_0__7__N_3441[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[173] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i663.GSR = "ENABLED";
    FD1P3AX array_255___i664 (.D(array_0__7__N_3441[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[173] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i664.GSR = "ENABLED";
    FD1P3AX array_255___i665 (.D(array_0__7__N_3433[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[172] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i665.GSR = "ENABLED";
    FD1P3AX array_255___i666 (.D(array_0__7__N_3433[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[172] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i666.GSR = "ENABLED";
    FD1P3AX array_255___i667 (.D(array_0__7__N_3433[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[172] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i667.GSR = "ENABLED";
    FD1P3AX array_255___i668 (.D(array_0__7__N_3433[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[172] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i668.GSR = "ENABLED";
    FD1P3AX array_255___i669 (.D(array_0__7__N_3433[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[172] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i669.GSR = "ENABLED";
    FD1P3AX array_255___i670 (.D(array_0__7__N_3433[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[172] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i670.GSR = "ENABLED";
    FD1P3AX array_255___i671 (.D(array_0__7__N_3433[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[172] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i671.GSR = "ENABLED";
    FD1P3AX array_255___i672 (.D(array_0__7__N_3433[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[172] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i672.GSR = "ENABLED";
    FD1P3AX array_255___i673 (.D(array_0__7__N_3425[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[171] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i673.GSR = "ENABLED";
    FD1P3AX array_255___i674 (.D(array_0__7__N_3425[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[171] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i674.GSR = "ENABLED";
    FD1P3AX array_255___i675 (.D(array_0__7__N_3425[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[171] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i675.GSR = "ENABLED";
    FD1P3AX array_255___i676 (.D(array_0__7__N_3425[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[171] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i676.GSR = "ENABLED";
    FD1P3AX array_255___i677 (.D(array_0__7__N_3425[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[171] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i677.GSR = "ENABLED";
    FD1P3AX array_255___i678 (.D(array_0__7__N_3425[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[171] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i678.GSR = "ENABLED";
    FD1P3AX array_255___i679 (.D(array_0__7__N_3425[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[171] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i679.GSR = "ENABLED";
    FD1P3AX array_255___i680 (.D(array_0__7__N_3425[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[171] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i680.GSR = "ENABLED";
    FD1P3AX array_255___i681 (.D(array_0__7__N_3417[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[170] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i681.GSR = "ENABLED";
    FD1P3AX array_255___i682 (.D(array_0__7__N_3417[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[170] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i682.GSR = "ENABLED";
    FD1P3AX array_255___i683 (.D(array_0__7__N_3417[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[170] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i683.GSR = "ENABLED";
    FD1P3AX array_255___i684 (.D(array_0__7__N_3417[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[170] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i684.GSR = "ENABLED";
    FD1P3AX array_255___i685 (.D(array_0__7__N_3417[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[170] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i685.GSR = "ENABLED";
    FD1P3AX array_255___i686 (.D(array_0__7__N_3417[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[170] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i686.GSR = "ENABLED";
    FD1P3AX array_255___i687 (.D(array_0__7__N_3417[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[170] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i687.GSR = "ENABLED";
    FD1P3AX array_255___i688 (.D(array_0__7__N_3417[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[170] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i688.GSR = "ENABLED";
    FD1P3AX array_255___i689 (.D(array_0__7__N_3409[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[169] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i689.GSR = "ENABLED";
    FD1P3AX array_255___i690 (.D(array_0__7__N_3409[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[169] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i690.GSR = "ENABLED";
    FD1P3AX array_255___i691 (.D(array_0__7__N_3409[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[169] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i691.GSR = "ENABLED";
    FD1P3AX array_255___i692 (.D(array_0__7__N_3409[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[169] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i692.GSR = "ENABLED";
    FD1P3AX array_255___i693 (.D(array_0__7__N_3409[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[169] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i693.GSR = "ENABLED";
    FD1P3AX array_255___i694 (.D(array_0__7__N_3409[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[169] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i694.GSR = "ENABLED";
    FD1P3AX array_255___i695 (.D(array_0__7__N_3409[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[169] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i695.GSR = "ENABLED";
    FD1P3AX array_255___i696 (.D(array_0__7__N_3409[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[169] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i696.GSR = "ENABLED";
    FD1P3AX array_255___i697 (.D(array_0__7__N_3401[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[168] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i697.GSR = "ENABLED";
    FD1P3AX array_255___i698 (.D(array_0__7__N_3401[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[168] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i698.GSR = "ENABLED";
    FD1P3AX array_255___i699 (.D(array_0__7__N_3401[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[168] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i699.GSR = "ENABLED";
    FD1P3AX array_255___i700 (.D(array_0__7__N_3401[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[168] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i700.GSR = "ENABLED";
    FD1P3AX array_255___i701 (.D(array_0__7__N_3401[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[168] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i701.GSR = "ENABLED";
    FD1P3AX array_255___i702 (.D(array_0__7__N_3401[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[168] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i702.GSR = "ENABLED";
    FD1P3AX array_255___i703 (.D(array_0__7__N_3401[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[168] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i703.GSR = "ENABLED";
    FD1P3AX array_255___i704 (.D(array_0__7__N_3401[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[168] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i704.GSR = "ENABLED";
    FD1P3AX array_255___i705 (.D(array_0__7__N_3393[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[167] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i705.GSR = "ENABLED";
    FD1P3AX array_255___i706 (.D(array_0__7__N_3393[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[167] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i706.GSR = "ENABLED";
    FD1P3AX array_255___i707 (.D(array_0__7__N_3393[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[167] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i707.GSR = "ENABLED";
    FD1P3AX array_255___i708 (.D(array_0__7__N_3393[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[167] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i708.GSR = "ENABLED";
    FD1P3AX array_255___i709 (.D(array_0__7__N_3393[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[167] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i709.GSR = "ENABLED";
    FD1P3AX array_255___i710 (.D(array_0__7__N_3393[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[167] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i710.GSR = "ENABLED";
    FD1P3AX array_255___i711 (.D(array_0__7__N_3393[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[167] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i711.GSR = "ENABLED";
    FD1P3AX array_255___i712 (.D(array_0__7__N_3393[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[167] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i712.GSR = "ENABLED";
    FD1P3AX array_255___i713 (.D(array_0__7__N_3385[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[166] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i713.GSR = "ENABLED";
    FD1P3AX array_255___i714 (.D(array_0__7__N_3385[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[166] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i714.GSR = "ENABLED";
    FD1P3AX array_255___i715 (.D(array_0__7__N_3385[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[166] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i715.GSR = "ENABLED";
    FD1P3AX array_255___i716 (.D(array_0__7__N_3385[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[166] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i716.GSR = "ENABLED";
    FD1P3AX array_255___i717 (.D(array_0__7__N_3385[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[166] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i717.GSR = "ENABLED";
    FD1P3AX array_255___i718 (.D(array_0__7__N_3385[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[166] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i718.GSR = "ENABLED";
    FD1P3AX array_255___i719 (.D(array_0__7__N_3385[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[166] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i719.GSR = "ENABLED";
    FD1P3AX array_255___i720 (.D(array_0__7__N_3385[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[166] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i720.GSR = "ENABLED";
    FD1P3AX array_255___i721 (.D(array_0__7__N_3377[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[165] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i721.GSR = "ENABLED";
    FD1P3AX array_255___i722 (.D(array_0__7__N_3377[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[165] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i722.GSR = "ENABLED";
    FD1P3AX array_255___i723 (.D(array_0__7__N_3377[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[165] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i723.GSR = "ENABLED";
    FD1P3AX array_255___i724 (.D(array_0__7__N_3377[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[165] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i724.GSR = "ENABLED";
    FD1P3AX array_255___i725 (.D(array_0__7__N_3377[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[165] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i725.GSR = "ENABLED";
    FD1P3AX array_255___i726 (.D(array_0__7__N_3377[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[165] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i726.GSR = "ENABLED";
    FD1P3AX array_255___i727 (.D(array_0__7__N_3377[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[165] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i727.GSR = "ENABLED";
    FD1P3AX array_255___i728 (.D(array_0__7__N_3377[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[165] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i728.GSR = "ENABLED";
    FD1P3AX array_255___i729 (.D(array_0__7__N_3369[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[164] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i729.GSR = "ENABLED";
    FD1P3AX array_255___i730 (.D(array_0__7__N_3369[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[164] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i730.GSR = "ENABLED";
    FD1P3AX array_255___i731 (.D(array_0__7__N_3369[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[164] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i731.GSR = "ENABLED";
    FD1P3AX array_255___i732 (.D(array_0__7__N_3369[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[164] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i732.GSR = "ENABLED";
    FD1P3AX array_255___i733 (.D(array_0__7__N_3369[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[164] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i733.GSR = "ENABLED";
    FD1P3AX array_255___i734 (.D(array_0__7__N_3369[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[164] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i734.GSR = "ENABLED";
    FD1P3AX array_255___i735 (.D(array_0__7__N_3369[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[164] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i735.GSR = "ENABLED";
    FD1P3AX array_255___i736 (.D(array_0__7__N_3369[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[164] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i736.GSR = "ENABLED";
    FD1P3AX array_255___i737 (.D(array_0__7__N_3361[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[163] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i737.GSR = "ENABLED";
    FD1P3AX array_255___i738 (.D(array_0__7__N_3361[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[163] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i738.GSR = "ENABLED";
    FD1P3AX array_255___i739 (.D(array_0__7__N_3361[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[163] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i739.GSR = "ENABLED";
    FD1P3AX array_255___i740 (.D(array_0__7__N_3361[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[163] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i740.GSR = "ENABLED";
    FD1P3AX array_255___i741 (.D(array_0__7__N_3361[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[163] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i741.GSR = "ENABLED";
    FD1P3AX array_255___i742 (.D(array_0__7__N_3361[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[163] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i742.GSR = "ENABLED";
    FD1P3AX array_255___i743 (.D(array_0__7__N_3361[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[163] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i743.GSR = "ENABLED";
    FD1P3AX array_255___i744 (.D(array_0__7__N_3361[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[163] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i744.GSR = "ENABLED";
    FD1P3AX array_255___i745 (.D(array_0__7__N_3353[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[162] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i745.GSR = "ENABLED";
    FD1P3AX array_255___i746 (.D(array_0__7__N_3353[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[162] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i746.GSR = "ENABLED";
    FD1P3AX array_255___i747 (.D(array_0__7__N_3353[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[162] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i747.GSR = "ENABLED";
    FD1P3AX array_255___i748 (.D(array_0__7__N_3353[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[162] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i748.GSR = "ENABLED";
    FD1P3AX array_255___i749 (.D(array_0__7__N_3353[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[162] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i749.GSR = "ENABLED";
    FD1P3AX array_255___i750 (.D(array_0__7__N_3353[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[162] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i750.GSR = "ENABLED";
    FD1P3AX array_255___i751 (.D(array_0__7__N_3353[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[162] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i751.GSR = "ENABLED";
    FD1P3AX array_255___i752 (.D(array_0__7__N_3353[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[162] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i752.GSR = "ENABLED";
    FD1P3AX array_255___i753 (.D(array_0__7__N_3345[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[161] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i753.GSR = "ENABLED";
    FD1P3AX array_255___i754 (.D(array_0__7__N_3345[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[161] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i754.GSR = "ENABLED";
    FD1P3AX array_255___i755 (.D(array_0__7__N_3345[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[161] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i755.GSR = "ENABLED";
    FD1P3AX array_255___i756 (.D(array_0__7__N_3345[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[161] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i756.GSR = "ENABLED";
    FD1P3AX array_255___i757 (.D(array_0__7__N_3345[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[161] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i757.GSR = "ENABLED";
    FD1P3AX array_255___i758 (.D(array_0__7__N_3345[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[161] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i758.GSR = "ENABLED";
    FD1P3AX array_255___i759 (.D(array_0__7__N_3345[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[161] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i759.GSR = "ENABLED";
    FD1P3AX array_255___i760 (.D(array_0__7__N_3345[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[161] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i760.GSR = "ENABLED";
    FD1P3AX array_255___i761 (.D(array_0__7__N_3337[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[160] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i761.GSR = "ENABLED";
    FD1P3AX array_255___i762 (.D(array_0__7__N_3337[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[160] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i762.GSR = "ENABLED";
    FD1P3AX array_255___i763 (.D(array_0__7__N_3337[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[160] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i763.GSR = "ENABLED";
    FD1P3AX array_255___i764 (.D(array_0__7__N_3337[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[160] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i764.GSR = "ENABLED";
    FD1P3AX array_255___i765 (.D(array_0__7__N_3337[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[160] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i765.GSR = "ENABLED";
    FD1P3AX array_255___i766 (.D(array_0__7__N_3337[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[160] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i766.GSR = "ENABLED";
    FD1P3AX array_255___i767 (.D(array_0__7__N_3337[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[160] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i767.GSR = "ENABLED";
    FD1P3AX array_255___i768 (.D(array_0__7__N_3337[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[160] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i768.GSR = "ENABLED";
    FD1P3AX array_255___i769 (.D(array_0__7__N_3329[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[159] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i769.GSR = "ENABLED";
    FD1P3AX array_255___i770 (.D(array_0__7__N_3329[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[159] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i770.GSR = "ENABLED";
    FD1P3AX array_255___i771 (.D(array_0__7__N_3329[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[159] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i771.GSR = "ENABLED";
    FD1P3AX array_255___i772 (.D(array_0__7__N_3329[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[159] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i772.GSR = "ENABLED";
    FD1P3AX array_255___i773 (.D(array_0__7__N_3329[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[159] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i773.GSR = "ENABLED";
    FD1P3AX array_255___i774 (.D(array_0__7__N_3329[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[159] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i774.GSR = "ENABLED";
    FD1P3AX array_255___i775 (.D(array_0__7__N_3329[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[159] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i775.GSR = "ENABLED";
    FD1P3AX array_255___i776 (.D(array_0__7__N_3329[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[159] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i776.GSR = "ENABLED";
    FD1P3AX array_255___i777 (.D(array_0__7__N_3321[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[158] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i777.GSR = "ENABLED";
    FD1P3AX array_255___i778 (.D(array_0__7__N_3321[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[158] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i778.GSR = "ENABLED";
    FD1P3AX array_255___i779 (.D(array_0__7__N_3321[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[158] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i779.GSR = "ENABLED";
    FD1P3AX array_255___i780 (.D(array_0__7__N_3321[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[158] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i780.GSR = "ENABLED";
    FD1P3AX array_255___i781 (.D(array_0__7__N_3321[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[158] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i781.GSR = "ENABLED";
    FD1P3AX array_255___i782 (.D(array_0__7__N_3321[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[158] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i782.GSR = "ENABLED";
    FD1P3AX array_255___i783 (.D(array_0__7__N_3321[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[158] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i783.GSR = "ENABLED";
    FD1P3AX array_255___i784 (.D(array_0__7__N_3321[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[158] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i784.GSR = "ENABLED";
    FD1P3AX array_255___i785 (.D(array_0__7__N_3313[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[157] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i785.GSR = "ENABLED";
    FD1P3AX array_255___i786 (.D(array_0__7__N_3313[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[157] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i786.GSR = "ENABLED";
    FD1P3AX array_255___i787 (.D(array_0__7__N_3313[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[157] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i787.GSR = "ENABLED";
    FD1P3AX array_255___i788 (.D(array_0__7__N_3313[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[157] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i788.GSR = "ENABLED";
    FD1P3AX array_255___i789 (.D(array_0__7__N_3313[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[157] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i789.GSR = "ENABLED";
    FD1P3AX array_255___i790 (.D(array_0__7__N_3313[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[157] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i790.GSR = "ENABLED";
    FD1P3AX array_255___i791 (.D(array_0__7__N_3313[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[157] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i791.GSR = "ENABLED";
    FD1P3AX array_255___i792 (.D(array_0__7__N_3313[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[157] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i792.GSR = "ENABLED";
    FD1P3AX array_255___i793 (.D(array_0__7__N_3305[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[156] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i793.GSR = "ENABLED";
    FD1P3AX array_255___i794 (.D(array_0__7__N_3305[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[156] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i794.GSR = "ENABLED";
    FD1P3AX array_255___i795 (.D(array_0__7__N_3305[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[156] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i795.GSR = "ENABLED";
    FD1P3AX array_255___i796 (.D(array_0__7__N_3305[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[156] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i796.GSR = "ENABLED";
    FD1P3AX array_255___i797 (.D(array_0__7__N_3305[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[156] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i797.GSR = "ENABLED";
    FD1P3AX array_255___i798 (.D(array_0__7__N_3305[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[156] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i798.GSR = "ENABLED";
    FD1P3AX array_255___i799 (.D(array_0__7__N_3305[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[156] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i799.GSR = "ENABLED";
    FD1P3AX array_255___i800 (.D(array_0__7__N_3305[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[156] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i800.GSR = "ENABLED";
    FD1P3AX array_255___i801 (.D(array_0__7__N_3297[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[155] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i801.GSR = "ENABLED";
    FD1P3AX array_255___i802 (.D(array_0__7__N_3297[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[155] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i802.GSR = "ENABLED";
    FD1P3AX array_255___i803 (.D(array_0__7__N_3297[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[155] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i803.GSR = "ENABLED";
    FD1P3AX array_255___i804 (.D(array_0__7__N_3297[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[155] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i804.GSR = "ENABLED";
    FD1P3AX array_255___i805 (.D(array_0__7__N_3297[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[155] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i805.GSR = "ENABLED";
    FD1P3AX array_255___i806 (.D(array_0__7__N_3297[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[155] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i806.GSR = "ENABLED";
    FD1P3AX array_255___i807 (.D(array_0__7__N_3297[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[155] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i807.GSR = "ENABLED";
    FD1P3AX array_255___i808 (.D(array_0__7__N_3297[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[155] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i808.GSR = "ENABLED";
    FD1P3AX array_255___i809 (.D(array_0__7__N_3289[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[154] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i809.GSR = "ENABLED";
    FD1P3AX array_255___i810 (.D(array_0__7__N_3289[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[154] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i810.GSR = "ENABLED";
    FD1P3AX array_255___i811 (.D(array_0__7__N_3289[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[154] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i811.GSR = "ENABLED";
    FD1P3AX array_255___i812 (.D(array_0__7__N_3289[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[154] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i812.GSR = "ENABLED";
    FD1P3AX array_255___i813 (.D(array_0__7__N_3289[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[154] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i813.GSR = "ENABLED";
    FD1P3AX array_255___i814 (.D(array_0__7__N_3289[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[154] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i814.GSR = "ENABLED";
    FD1P3AX array_255___i815 (.D(array_0__7__N_3289[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[154] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i815.GSR = "ENABLED";
    FD1P3AX array_255___i816 (.D(array_0__7__N_3289[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[154] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i816.GSR = "ENABLED";
    FD1P3AX array_255___i817 (.D(array_0__7__N_3281[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[153] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i817.GSR = "ENABLED";
    FD1P3AX array_255___i818 (.D(array_0__7__N_3281[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[153] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i818.GSR = "ENABLED";
    FD1P3AX array_255___i819 (.D(array_0__7__N_3281[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[153] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i819.GSR = "ENABLED";
    FD1P3AX array_255___i820 (.D(array_0__7__N_3281[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[153] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i820.GSR = "ENABLED";
    FD1P3AX array_255___i821 (.D(array_0__7__N_3281[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[153] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i821.GSR = "ENABLED";
    FD1P3AX array_255___i822 (.D(array_0__7__N_3281[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[153] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i822.GSR = "ENABLED";
    FD1P3AX array_255___i823 (.D(array_0__7__N_3281[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[153] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i823.GSR = "ENABLED";
    FD1P3AX array_255___i824 (.D(array_0__7__N_3281[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[153] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i824.GSR = "ENABLED";
    FD1P3AX array_255___i825 (.D(array_0__7__N_3273[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[152] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i825.GSR = "ENABLED";
    FD1P3AX array_255___i826 (.D(array_0__7__N_3273[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[152] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i826.GSR = "ENABLED";
    FD1P3AX array_255___i827 (.D(array_0__7__N_3273[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[152] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i827.GSR = "ENABLED";
    FD1P3AX array_255___i828 (.D(array_0__7__N_3273[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[152] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i828.GSR = "ENABLED";
    FD1P3AX array_255___i829 (.D(array_0__7__N_3273[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[152] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i829.GSR = "ENABLED";
    FD1P3AX array_255___i830 (.D(array_0__7__N_3273[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[152] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i830.GSR = "ENABLED";
    FD1P3AX array_255___i831 (.D(array_0__7__N_3273[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[152] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i831.GSR = "ENABLED";
    FD1P3AX array_255___i832 (.D(array_0__7__N_3273[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[152] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i832.GSR = "ENABLED";
    FD1P3AX array_255___i833 (.D(array_0__7__N_3265[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[151] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i833.GSR = "ENABLED";
    FD1P3AX array_255___i834 (.D(array_0__7__N_3265[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[151] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i834.GSR = "ENABLED";
    FD1P3AX array_255___i835 (.D(array_0__7__N_3265[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[151] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i835.GSR = "ENABLED";
    FD1P3AX array_255___i836 (.D(array_0__7__N_3265[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[151] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i836.GSR = "ENABLED";
    FD1P3AX array_255___i837 (.D(array_0__7__N_3265[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[151] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i837.GSR = "ENABLED";
    FD1P3AX array_255___i838 (.D(array_0__7__N_3265[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[151] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i838.GSR = "ENABLED";
    FD1P3AX array_255___i839 (.D(array_0__7__N_3265[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[151] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i839.GSR = "ENABLED";
    FD1P3AX array_255___i840 (.D(array_0__7__N_3265[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[151] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i840.GSR = "ENABLED";
    FD1P3AX array_255___i841 (.D(array_0__7__N_3257[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[150] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i841.GSR = "ENABLED";
    FD1P3AX array_255___i842 (.D(array_0__7__N_3257[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[150] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i842.GSR = "ENABLED";
    FD1P3AX array_255___i843 (.D(array_0__7__N_3257[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[150] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i843.GSR = "ENABLED";
    FD1P3AX array_255___i844 (.D(array_0__7__N_3257[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[150] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i844.GSR = "ENABLED";
    FD1P3AX array_255___i845 (.D(array_0__7__N_3257[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[150] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i845.GSR = "ENABLED";
    FD1P3AX array_255___i846 (.D(array_0__7__N_3257[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[150] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i846.GSR = "ENABLED";
    FD1P3AX array_255___i847 (.D(array_0__7__N_3257[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[150] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i847.GSR = "ENABLED";
    FD1P3AX array_255___i848 (.D(array_0__7__N_3257[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[150] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i848.GSR = "ENABLED";
    FD1P3AX array_255___i849 (.D(array_0__7__N_3249[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[149] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i849.GSR = "ENABLED";
    FD1P3AX array_255___i850 (.D(array_0__7__N_3249[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[149] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i850.GSR = "ENABLED";
    FD1P3AX array_255___i851 (.D(array_0__7__N_3249[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[149] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i851.GSR = "ENABLED";
    FD1P3AX array_255___i852 (.D(array_0__7__N_3249[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[149] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i852.GSR = "ENABLED";
    FD1P3AX array_255___i853 (.D(array_0__7__N_3249[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[149] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i853.GSR = "ENABLED";
    FD1P3AX array_255___i854 (.D(array_0__7__N_3249[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[149] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i854.GSR = "ENABLED";
    FD1P3AX array_255___i855 (.D(array_0__7__N_3249[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[149] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i855.GSR = "ENABLED";
    FD1P3AX array_255___i856 (.D(array_0__7__N_3249[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[149] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i856.GSR = "ENABLED";
    FD1P3AX array_255___i857 (.D(array_0__7__N_3241[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[148] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i857.GSR = "ENABLED";
    FD1P3AX array_255___i858 (.D(array_0__7__N_3241[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[148] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i858.GSR = "ENABLED";
    FD1P3AX array_255___i859 (.D(array_0__7__N_3241[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[148] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i859.GSR = "ENABLED";
    FD1P3AX array_255___i860 (.D(array_0__7__N_3241[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[148] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i860.GSR = "ENABLED";
    FD1P3AX array_255___i861 (.D(array_0__7__N_3241[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[148] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i861.GSR = "ENABLED";
    FD1P3AX array_255___i862 (.D(array_0__7__N_3241[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[148] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i862.GSR = "ENABLED";
    FD1P3AX array_255___i863 (.D(array_0__7__N_3241[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[148] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i863.GSR = "ENABLED";
    FD1P3AX array_255___i864 (.D(array_0__7__N_3241[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[148] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i864.GSR = "ENABLED";
    FD1P3AX array_255___i865 (.D(array_0__7__N_3233[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[147] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i865.GSR = "ENABLED";
    FD1P3AX array_255___i866 (.D(array_0__7__N_3233[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[147] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i866.GSR = "ENABLED";
    FD1P3AX array_255___i867 (.D(array_0__7__N_3233[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[147] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i867.GSR = "ENABLED";
    FD1P3AX array_255___i868 (.D(array_0__7__N_3233[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[147] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i868.GSR = "ENABLED";
    FD1P3AX array_255___i869 (.D(array_0__7__N_3233[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[147] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i869.GSR = "ENABLED";
    FD1P3AX array_255___i870 (.D(array_0__7__N_3233[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[147] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i870.GSR = "ENABLED";
    FD1P3AX array_255___i871 (.D(array_0__7__N_3233[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[147] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i871.GSR = "ENABLED";
    FD1P3AX array_255___i872 (.D(array_0__7__N_3233[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[147] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i872.GSR = "ENABLED";
    FD1P3AX array_255___i873 (.D(array_0__7__N_3225[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[146] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i873.GSR = "ENABLED";
    FD1P3AX array_255___i874 (.D(array_0__7__N_3225[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[146] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i874.GSR = "ENABLED";
    FD1P3AX array_255___i875 (.D(array_0__7__N_3225[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[146] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i875.GSR = "ENABLED";
    FD1P3AX array_255___i876 (.D(array_0__7__N_3225[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[146] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i876.GSR = "ENABLED";
    FD1P3AX array_255___i877 (.D(array_0__7__N_3225[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[146] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i877.GSR = "ENABLED";
    FD1P3AX array_255___i878 (.D(array_0__7__N_3225[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[146] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i878.GSR = "ENABLED";
    FD1P3AX array_255___i879 (.D(array_0__7__N_3225[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[146] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i879.GSR = "ENABLED";
    FD1P3AX array_255___i880 (.D(array_0__7__N_3225[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[146] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i880.GSR = "ENABLED";
    FD1P3AX array_255___i881 (.D(array_0__7__N_3217[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[145] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i881.GSR = "ENABLED";
    FD1P3AX array_255___i882 (.D(array_0__7__N_3217[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[145] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i882.GSR = "ENABLED";
    FD1P3AX array_255___i883 (.D(array_0__7__N_3217[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[145] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i883.GSR = "ENABLED";
    FD1P3AX array_255___i884 (.D(array_0__7__N_3217[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[145] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i884.GSR = "ENABLED";
    FD1P3AX array_255___i885 (.D(array_0__7__N_3217[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[145] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i885.GSR = "ENABLED";
    FD1P3AX array_255___i886 (.D(array_0__7__N_3217[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[145] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i886.GSR = "ENABLED";
    FD1P3AX array_255___i887 (.D(array_0__7__N_3217[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[145] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i887.GSR = "ENABLED";
    FD1P3AX array_255___i888 (.D(array_0__7__N_3217[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[145] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i888.GSR = "ENABLED";
    FD1P3AX array_255___i889 (.D(array_0__7__N_3209[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[144] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i889.GSR = "ENABLED";
    FD1P3AX array_255___i890 (.D(array_0__7__N_3209[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[144] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i890.GSR = "ENABLED";
    FD1P3AX array_255___i891 (.D(array_0__7__N_3209[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[144] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i891.GSR = "ENABLED";
    FD1P3AX array_255___i892 (.D(array_0__7__N_3209[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[144] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i892.GSR = "ENABLED";
    FD1P3AX array_255___i893 (.D(array_0__7__N_3209[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[144] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i893.GSR = "ENABLED";
    FD1P3AX array_255___i894 (.D(array_0__7__N_3209[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[144] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i894.GSR = "ENABLED";
    FD1P3AX array_255___i895 (.D(array_0__7__N_3209[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[144] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i895.GSR = "ENABLED";
    FD1P3AX array_255___i896 (.D(array_0__7__N_3209[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[144] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i896.GSR = "ENABLED";
    FD1P3AX array_255___i897 (.D(array_0__7__N_3201[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[143] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i897.GSR = "ENABLED";
    FD1P3AX array_255___i898 (.D(array_0__7__N_3201[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[143] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i898.GSR = "ENABLED";
    FD1P3AX array_255___i899 (.D(array_0__7__N_3201[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[143] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i899.GSR = "ENABLED";
    FD1P3AX array_255___i900 (.D(array_0__7__N_3201[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[143] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i900.GSR = "ENABLED";
    FD1P3AX array_255___i901 (.D(array_0__7__N_3201[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[143] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i901.GSR = "ENABLED";
    FD1P3AX array_255___i902 (.D(array_0__7__N_3201[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[143] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i902.GSR = "ENABLED";
    FD1P3AX array_255___i903 (.D(array_0__7__N_3201[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[143] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i903.GSR = "ENABLED";
    FD1P3AX array_255___i904 (.D(array_0__7__N_3201[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[143] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i904.GSR = "ENABLED";
    FD1P3AX array_255___i905 (.D(array_0__7__N_3193[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[142] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i905.GSR = "ENABLED";
    FD1P3AX array_255___i906 (.D(array_0__7__N_3193[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[142] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i906.GSR = "ENABLED";
    FD1P3AX array_255___i907 (.D(array_0__7__N_3193[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[142] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i907.GSR = "ENABLED";
    FD1P3AX array_255___i908 (.D(array_0__7__N_3193[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[142] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i908.GSR = "ENABLED";
    FD1P3AX array_255___i909 (.D(array_0__7__N_3193[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[142] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i909.GSR = "ENABLED";
    FD1P3AX array_255___i910 (.D(array_0__7__N_3193[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[142] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i910.GSR = "ENABLED";
    FD1P3AX array_255___i911 (.D(array_0__7__N_3193[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[142] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i911.GSR = "ENABLED";
    FD1P3AX array_255___i912 (.D(array_0__7__N_3193[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[142] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i912.GSR = "ENABLED";
    FD1P3AX array_255___i913 (.D(array_0__7__N_3185[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[141] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i913.GSR = "ENABLED";
    FD1P3AX array_255___i914 (.D(array_0__7__N_3185[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[141] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i914.GSR = "ENABLED";
    FD1P3AX array_255___i915 (.D(array_0__7__N_3185[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[141] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i915.GSR = "ENABLED";
    FD1P3AX array_255___i916 (.D(array_0__7__N_3185[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[141] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i916.GSR = "ENABLED";
    FD1P3AX array_255___i917 (.D(array_0__7__N_3185[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[141] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i917.GSR = "ENABLED";
    FD1P3AX array_255___i918 (.D(array_0__7__N_3185[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[141] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i918.GSR = "ENABLED";
    FD1P3AX array_255___i919 (.D(array_0__7__N_3185[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[141] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i919.GSR = "ENABLED";
    FD1P3AX array_255___i920 (.D(array_0__7__N_3185[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[141] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i920.GSR = "ENABLED";
    FD1P3AX array_255___i921 (.D(array_0__7__N_3177[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[140] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i921.GSR = "ENABLED";
    FD1P3AX array_255___i922 (.D(array_0__7__N_3177[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[140] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i922.GSR = "ENABLED";
    FD1P3AX array_255___i923 (.D(array_0__7__N_3177[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[140] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i923.GSR = "ENABLED";
    FD1P3AX array_255___i924 (.D(array_0__7__N_3177[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[140] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i924.GSR = "ENABLED";
    FD1P3AX array_255___i925 (.D(array_0__7__N_3177[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[140] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i925.GSR = "ENABLED";
    FD1P3AX array_255___i926 (.D(array_0__7__N_3177[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[140] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i926.GSR = "ENABLED";
    FD1P3AX array_255___i927 (.D(array_0__7__N_3177[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[140] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i927.GSR = "ENABLED";
    FD1P3AX array_255___i928 (.D(array_0__7__N_3177[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[140] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i928.GSR = "ENABLED";
    FD1P3AX array_255___i929 (.D(array_0__7__N_3169[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[139] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i929.GSR = "ENABLED";
    FD1P3AX array_255___i930 (.D(array_0__7__N_3169[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[139] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i930.GSR = "ENABLED";
    FD1P3AX array_255___i931 (.D(array_0__7__N_3169[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[139] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i931.GSR = "ENABLED";
    FD1P3AX array_255___i932 (.D(array_0__7__N_3169[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[139] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i932.GSR = "ENABLED";
    FD1P3AX array_255___i933 (.D(array_0__7__N_3169[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[139] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i933.GSR = "ENABLED";
    FD1P3AX array_255___i934 (.D(array_0__7__N_3169[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[139] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i934.GSR = "ENABLED";
    FD1P3AX array_255___i935 (.D(array_0__7__N_3169[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[139] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i935.GSR = "ENABLED";
    FD1P3AX array_255___i936 (.D(array_0__7__N_3169[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[139] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i936.GSR = "ENABLED";
    FD1P3AX array_255___i937 (.D(array_0__7__N_3161[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[138] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i937.GSR = "ENABLED";
    FD1P3AX array_255___i938 (.D(array_0__7__N_3161[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[138] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i938.GSR = "ENABLED";
    FD1P3AX array_255___i939 (.D(array_0__7__N_3161[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[138] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i939.GSR = "ENABLED";
    FD1P3AX array_255___i940 (.D(array_0__7__N_3161[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[138] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i940.GSR = "ENABLED";
    FD1P3AX array_255___i941 (.D(array_0__7__N_3161[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[138] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i941.GSR = "ENABLED";
    FD1P3AX array_255___i942 (.D(array_0__7__N_3161[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[138] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i942.GSR = "ENABLED";
    FD1P3AX array_255___i943 (.D(array_0__7__N_3161[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[138] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i943.GSR = "ENABLED";
    FD1P3AX array_255___i944 (.D(array_0__7__N_3161[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[138] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i944.GSR = "ENABLED";
    FD1P3AX array_255___i945 (.D(array_0__7__N_3153[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[137] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i945.GSR = "ENABLED";
    FD1P3AX array_255___i946 (.D(array_0__7__N_3153[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[137] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i946.GSR = "ENABLED";
    FD1P3AX array_255___i947 (.D(array_0__7__N_3153[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[137] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i947.GSR = "ENABLED";
    FD1P3AX array_255___i948 (.D(array_0__7__N_3153[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[137] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i948.GSR = "ENABLED";
    FD1P3AX array_255___i949 (.D(array_0__7__N_3153[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[137] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i949.GSR = "ENABLED";
    FD1P3AX array_255___i950 (.D(array_0__7__N_3153[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[137] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i950.GSR = "ENABLED";
    FD1P3AX array_255___i951 (.D(array_0__7__N_3153[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[137] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i951.GSR = "ENABLED";
    FD1P3AX array_255___i952 (.D(array_0__7__N_3153[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[137] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i952.GSR = "ENABLED";
    FD1P3AX array_255___i953 (.D(array_0__7__N_3145[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[136] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i953.GSR = "ENABLED";
    FD1P3AX array_255___i954 (.D(array_0__7__N_3145[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[136] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i954.GSR = "ENABLED";
    FD1P3AX array_255___i955 (.D(array_0__7__N_3145[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[136] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i955.GSR = "ENABLED";
    FD1P3AX array_255___i956 (.D(array_0__7__N_3145[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[136] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i956.GSR = "ENABLED";
    FD1P3AX array_255___i957 (.D(array_0__7__N_3145[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[136] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i957.GSR = "ENABLED";
    FD1P3AX array_255___i958 (.D(array_0__7__N_3145[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[136] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i958.GSR = "ENABLED";
    FD1P3AX array_255___i959 (.D(array_0__7__N_3145[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[136] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i959.GSR = "ENABLED";
    FD1P3AX array_255___i960 (.D(array_0__7__N_3145[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[136] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i960.GSR = "ENABLED";
    FD1P3AX array_255___i961 (.D(array_0__7__N_3137[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[135] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i961.GSR = "ENABLED";
    FD1P3AX array_255___i962 (.D(array_0__7__N_3137[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[135] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i962.GSR = "ENABLED";
    FD1P3AX array_255___i963 (.D(array_0__7__N_3137[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[135] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i963.GSR = "ENABLED";
    FD1P3AX array_255___i964 (.D(array_0__7__N_3137[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[135] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i964.GSR = "ENABLED";
    FD1P3AX array_255___i965 (.D(array_0__7__N_3137[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[135] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i965.GSR = "ENABLED";
    FD1P3AX array_255___i966 (.D(array_0__7__N_3137[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[135] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i966.GSR = "ENABLED";
    FD1P3AX array_255___i967 (.D(array_0__7__N_3137[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[135] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i967.GSR = "ENABLED";
    FD1P3AX array_255___i968 (.D(array_0__7__N_3137[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[135] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i968.GSR = "ENABLED";
    FD1P3AX array_255___i969 (.D(array_0__7__N_3129[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[134] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i969.GSR = "ENABLED";
    FD1P3AX array_255___i970 (.D(array_0__7__N_3129[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[134] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i970.GSR = "ENABLED";
    FD1P3AX array_255___i971 (.D(array_0__7__N_3129[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[134] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i971.GSR = "ENABLED";
    FD1P3AX array_255___i972 (.D(array_0__7__N_3129[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[134] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i972.GSR = "ENABLED";
    FD1P3AX array_255___i973 (.D(array_0__7__N_3129[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[134] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i973.GSR = "ENABLED";
    FD1P3AX array_255___i974 (.D(array_0__7__N_3129[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[134] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i974.GSR = "ENABLED";
    FD1P3AX array_255___i975 (.D(array_0__7__N_3129[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[134] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i975.GSR = "ENABLED";
    FD1P3AX array_255___i976 (.D(array_0__7__N_3129[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[134] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i976.GSR = "ENABLED";
    FD1P3AX array_255___i977 (.D(array_0__7__N_3121[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[133] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i977.GSR = "ENABLED";
    FD1P3AX array_255___i978 (.D(array_0__7__N_3121[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[133] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i978.GSR = "ENABLED";
    FD1P3AX array_255___i979 (.D(array_0__7__N_3121[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[133] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i979.GSR = "ENABLED";
    FD1P3AX array_255___i980 (.D(array_0__7__N_3121[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[133] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i980.GSR = "ENABLED";
    FD1P3AX array_255___i981 (.D(array_0__7__N_3121[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[133] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i981.GSR = "ENABLED";
    FD1P3AX array_255___i982 (.D(array_0__7__N_3121[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[133] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i982.GSR = "ENABLED";
    FD1P3AX array_255___i983 (.D(array_0__7__N_3121[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[133] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i983.GSR = "ENABLED";
    FD1P3AX array_255___i984 (.D(array_0__7__N_3121[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[133] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i984.GSR = "ENABLED";
    FD1P3AX array_255___i985 (.D(array_0__7__N_3113[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[132] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i985.GSR = "ENABLED";
    FD1P3AX array_255___i986 (.D(array_0__7__N_3113[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[132] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i986.GSR = "ENABLED";
    FD1P3AX array_255___i987 (.D(array_0__7__N_3113[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[132] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i987.GSR = "ENABLED";
    FD1P3AX array_255___i988 (.D(array_0__7__N_3113[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[132] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i988.GSR = "ENABLED";
    FD1P3AX array_255___i989 (.D(array_0__7__N_3113[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[132] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i989.GSR = "ENABLED";
    FD1P3AX array_255___i990 (.D(array_0__7__N_3113[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[132] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i990.GSR = "ENABLED";
    FD1P3AX array_255___i991 (.D(array_0__7__N_3113[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[132] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i991.GSR = "ENABLED";
    FD1P3AX array_255___i992 (.D(array_0__7__N_3113[7]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[132] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i992.GSR = "ENABLED";
    FD1P3AX array_255___i993 (.D(array_0__7__N_3105[0]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[131] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i993.GSR = "ENABLED";
    FD1P3AX array_255___i994 (.D(array_0__7__N_3105[1]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[131] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i994.GSR = "ENABLED";
    FD1P3AX array_255___i995 (.D(array_0__7__N_3105[2]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[131] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i995.GSR = "ENABLED";
    FD1P3AX array_255___i996 (.D(array_0__7__N_3105[3]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[131] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i996.GSR = "ENABLED";
    FD1P3AX array_255___i997 (.D(array_0__7__N_3105[4]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[131] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i997.GSR = "ENABLED";
    FD1P3AX array_255___i998 (.D(array_0__7__N_3105[5]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[131] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i998.GSR = "ENABLED";
    FD1P3AX array_255___i999 (.D(array_0__7__N_3105[6]), .SP(clk_c_enable_1007), 
            .CK(clk_c), .Q(\array[131] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i999.GSR = "ENABLED";
    FD1P3AX array_255___i1000 (.D(array_0__7__N_3105[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[131] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1000.GSR = "ENABLED";
    FD1P3AX array_255___i1001 (.D(array_0__7__N_3097[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[130] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1001.GSR = "ENABLED";
    FD1P3AX array_255___i1002 (.D(array_0__7__N_3097[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[130] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1002.GSR = "ENABLED";
    FD1P3AX array_255___i1003 (.D(array_0__7__N_3097[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[130] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1003.GSR = "ENABLED";
    FD1P3AX array_255___i1004 (.D(array_0__7__N_3097[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[130] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1004.GSR = "ENABLED";
    FD1P3AX array_255___i1005 (.D(array_0__7__N_3097[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[130] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1005.GSR = "ENABLED";
    FD1P3AX array_255___i1006 (.D(array_0__7__N_3097[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[130] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1006.GSR = "ENABLED";
    FD1P3AX array_255___i1007 (.D(array_0__7__N_3097[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[130] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1007.GSR = "ENABLED";
    FD1P3AX array_255___i1008 (.D(array_0__7__N_3097[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[130] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1008.GSR = "ENABLED";
    FD1P3AX array_255___i1009 (.D(array_0__7__N_3089[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[129] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1009.GSR = "ENABLED";
    FD1P3AX array_255___i1010 (.D(array_0__7__N_3089[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[129] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1010.GSR = "ENABLED";
    FD1P3AX array_255___i1011 (.D(array_0__7__N_3089[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[129] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1011.GSR = "ENABLED";
    FD1P3AX array_255___i1012 (.D(array_0__7__N_3089[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[129] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1012.GSR = "ENABLED";
    FD1P3AX array_255___i1013 (.D(array_0__7__N_3089[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[129] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1013.GSR = "ENABLED";
    FD1P3AX array_255___i1014 (.D(array_0__7__N_3089[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[129] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1014.GSR = "ENABLED";
    FD1P3AX array_255___i1015 (.D(array_0__7__N_3089[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[129] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1015.GSR = "ENABLED";
    FD1P3AX array_255___i1016 (.D(array_0__7__N_3089[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[129] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1016.GSR = "ENABLED";
    FD1P3AX array_255___i1017 (.D(array_0__7__N_3081[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[128] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1017.GSR = "ENABLED";
    FD1P3AX array_255___i1018 (.D(array_0__7__N_3081[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[128] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1018.GSR = "ENABLED";
    FD1P3AX array_255___i1019 (.D(array_0__7__N_3081[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[128] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1019.GSR = "ENABLED";
    FD1P3AX array_255___i1020 (.D(array_0__7__N_3081[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[128] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1020.GSR = "ENABLED";
    FD1P3AX array_255___i1021 (.D(array_0__7__N_3081[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[128] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1021.GSR = "ENABLED";
    FD1P3AX array_255___i1022 (.D(array_0__7__N_3081[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[128] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1022.GSR = "ENABLED";
    FD1P3AX array_255___i1023 (.D(array_0__7__N_3081[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[128] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1023.GSR = "ENABLED";
    FD1P3AX array_255___i1024 (.D(array_0__7__N_3081[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[128] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1024.GSR = "ENABLED";
    FD1P3AX array_255___i1025 (.D(array_0__7__N_3073[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[127] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1025.GSR = "ENABLED";
    FD1P3AX array_255___i1026 (.D(array_0__7__N_3073[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[127] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1026.GSR = "ENABLED";
    FD1P3AX array_255___i1027 (.D(array_0__7__N_3073[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[127] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1027.GSR = "ENABLED";
    FD1P3AX array_255___i1028 (.D(array_0__7__N_3073[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[127] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1028.GSR = "ENABLED";
    FD1P3AX array_255___i1029 (.D(array_0__7__N_3073[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[127] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1029.GSR = "ENABLED";
    FD1P3AX array_255___i1030 (.D(array_0__7__N_3073[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[127] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1030.GSR = "ENABLED";
    FD1P3AX array_255___i1031 (.D(array_0__7__N_3073[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[127] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1031.GSR = "ENABLED";
    FD1P3AX array_255___i1032 (.D(array_0__7__N_3073[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[127] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1032.GSR = "ENABLED";
    FD1P3AX array_255___i1033 (.D(array_0__7__N_3065[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[126] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1033.GSR = "ENABLED";
    FD1P3AX array_255___i1034 (.D(array_0__7__N_3065[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[126] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1034.GSR = "ENABLED";
    FD1P3AX array_255___i1035 (.D(array_0__7__N_3065[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[126] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1035.GSR = "ENABLED";
    FD1P3AX array_255___i1036 (.D(array_0__7__N_3065[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[126] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1036.GSR = "ENABLED";
    FD1P3AX array_255___i1037 (.D(array_0__7__N_3065[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[126] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1037.GSR = "ENABLED";
    FD1P3AX array_255___i1038 (.D(array_0__7__N_3065[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[126] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1038.GSR = "ENABLED";
    FD1P3AX array_255___i1039 (.D(array_0__7__N_3065[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[126] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1039.GSR = "ENABLED";
    FD1P3AX array_255___i1040 (.D(array_0__7__N_3065[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[126] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1040.GSR = "ENABLED";
    FD1P3AX array_255___i1041 (.D(array_0__7__N_3057[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[125] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1041.GSR = "ENABLED";
    FD1P3AX array_255___i1042 (.D(array_0__7__N_3057[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[125] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1042.GSR = "ENABLED";
    FD1P3AX array_255___i1043 (.D(array_0__7__N_3057[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[125] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1043.GSR = "ENABLED";
    FD1P3AX array_255___i1044 (.D(array_0__7__N_3057[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[125] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1044.GSR = "ENABLED";
    FD1P3AX array_255___i1045 (.D(array_0__7__N_3057[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[125] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1045.GSR = "ENABLED";
    FD1P3AX array_255___i1046 (.D(array_0__7__N_3057[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[125] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1046.GSR = "ENABLED";
    FD1P3AX array_255___i1047 (.D(array_0__7__N_3057[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[125] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1047.GSR = "ENABLED";
    FD1P3AX array_255___i1048 (.D(array_0__7__N_3057[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[125] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1048.GSR = "ENABLED";
    FD1P3AX array_255___i1049 (.D(array_0__7__N_3049[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[124] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1049.GSR = "ENABLED";
    FD1P3AX array_255___i1050 (.D(array_0__7__N_3049[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[124] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1050.GSR = "ENABLED";
    FD1P3AX array_255___i1051 (.D(array_0__7__N_3049[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[124] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1051.GSR = "ENABLED";
    FD1P3AX array_255___i1052 (.D(array_0__7__N_3049[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[124] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1052.GSR = "ENABLED";
    FD1P3AX array_255___i1053 (.D(array_0__7__N_3049[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[124] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1053.GSR = "ENABLED";
    FD1P3AX array_255___i1054 (.D(array_0__7__N_3049[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[124] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1054.GSR = "ENABLED";
    FD1P3AX array_255___i1055 (.D(array_0__7__N_3049[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[124] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1055.GSR = "ENABLED";
    FD1P3AX array_255___i1056 (.D(array_0__7__N_3049[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[124] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1056.GSR = "ENABLED";
    FD1P3AX array_255___i1057 (.D(array_0__7__N_3041[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[123] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1057.GSR = "ENABLED";
    FD1P3AX array_255___i1058 (.D(array_0__7__N_3041[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[123] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1058.GSR = "ENABLED";
    FD1P3AX array_255___i1059 (.D(array_0__7__N_3041[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[123] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1059.GSR = "ENABLED";
    FD1P3AX array_255___i1060 (.D(array_0__7__N_3041[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[123] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1060.GSR = "ENABLED";
    FD1P3AX array_255___i1061 (.D(array_0__7__N_3041[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[123] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1061.GSR = "ENABLED";
    FD1P3AX array_255___i1062 (.D(array_0__7__N_3041[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[123] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1062.GSR = "ENABLED";
    FD1P3AX array_255___i1063 (.D(array_0__7__N_3041[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[123] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1063.GSR = "ENABLED";
    FD1P3AX array_255___i1064 (.D(array_0__7__N_3041[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[123] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1064.GSR = "ENABLED";
    FD1P3AX array_255___i1065 (.D(array_0__7__N_3033[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[122] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1065.GSR = "ENABLED";
    FD1P3AX array_255___i1066 (.D(array_0__7__N_3033[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[122] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1066.GSR = "ENABLED";
    FD1P3AX array_255___i1067 (.D(array_0__7__N_3033[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[122] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1067.GSR = "ENABLED";
    FD1P3AX array_255___i1068 (.D(array_0__7__N_3033[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[122] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1068.GSR = "ENABLED";
    FD1P3AX array_255___i1069 (.D(array_0__7__N_3033[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[122] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1069.GSR = "ENABLED";
    FD1P3AX array_255___i1070 (.D(array_0__7__N_3033[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[122] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1070.GSR = "ENABLED";
    FD1P3AX array_255___i1071 (.D(array_0__7__N_3033[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[122] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1071.GSR = "ENABLED";
    FD1P3AX array_255___i1072 (.D(array_0__7__N_3033[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[122] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1072.GSR = "ENABLED";
    FD1P3AX array_255___i1073 (.D(array_0__7__N_3025[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[121] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1073.GSR = "ENABLED";
    FD1P3AX array_255___i1074 (.D(array_0__7__N_3025[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[121] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1074.GSR = "ENABLED";
    FD1P3AX array_255___i1075 (.D(array_0__7__N_3025[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[121] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1075.GSR = "ENABLED";
    FD1P3AX array_255___i1076 (.D(array_0__7__N_3025[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[121] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1076.GSR = "ENABLED";
    FD1P3AX array_255___i1077 (.D(array_0__7__N_3025[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[121] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1077.GSR = "ENABLED";
    FD1P3AX array_255___i1078 (.D(array_0__7__N_3025[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[121] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1078.GSR = "ENABLED";
    FD1P3AX array_255___i1079 (.D(array_0__7__N_3025[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[121] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1079.GSR = "ENABLED";
    FD1P3AX array_255___i1080 (.D(array_0__7__N_3025[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[121] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1080.GSR = "ENABLED";
    FD1P3AX array_255___i1081 (.D(array_0__7__N_3017[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[120] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1081.GSR = "ENABLED";
    FD1P3AX array_255___i1082 (.D(array_0__7__N_3017[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[120] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1082.GSR = "ENABLED";
    FD1P3AX array_255___i1083 (.D(array_0__7__N_3017[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[120] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1083.GSR = "ENABLED";
    FD1P3AX array_255___i1084 (.D(array_0__7__N_3017[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[120] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1084.GSR = "ENABLED";
    FD1P3AX array_255___i1085 (.D(array_0__7__N_3017[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[120] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1085.GSR = "ENABLED";
    FD1P3AX array_255___i1086 (.D(array_0__7__N_3017[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[120] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1086.GSR = "ENABLED";
    FD1P3AX array_255___i1087 (.D(array_0__7__N_3017[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[120] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1087.GSR = "ENABLED";
    FD1P3AX array_255___i1088 (.D(array_0__7__N_3017[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[120] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1088.GSR = "ENABLED";
    FD1P3AX array_255___i1089 (.D(array_0__7__N_3009[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[119] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1089.GSR = "ENABLED";
    FD1P3AX array_255___i1090 (.D(array_0__7__N_3009[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[119] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1090.GSR = "ENABLED";
    FD1P3AX array_255___i1091 (.D(array_0__7__N_3009[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[119] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1091.GSR = "ENABLED";
    FD1P3AX array_255___i1092 (.D(array_0__7__N_3009[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[119] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1092.GSR = "ENABLED";
    FD1P3AX array_255___i1093 (.D(array_0__7__N_3009[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[119] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1093.GSR = "ENABLED";
    FD1P3AX array_255___i1094 (.D(array_0__7__N_3009[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[119] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1094.GSR = "ENABLED";
    FD1P3AX array_255___i1095 (.D(array_0__7__N_3009[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[119] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1095.GSR = "ENABLED";
    FD1P3AX array_255___i1096 (.D(array_0__7__N_3009[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[119] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1096.GSR = "ENABLED";
    FD1P3AX array_255___i1097 (.D(array_0__7__N_3001[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[118] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1097.GSR = "ENABLED";
    FD1P3AX array_255___i1098 (.D(array_0__7__N_3001[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[118] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1098.GSR = "ENABLED";
    FD1P3AX array_255___i1099 (.D(array_0__7__N_3001[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[118] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1099.GSR = "ENABLED";
    FD1P3AX array_255___i1100 (.D(array_0__7__N_3001[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[118] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1100.GSR = "ENABLED";
    FD1P3AX array_255___i1101 (.D(array_0__7__N_3001[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[118] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1101.GSR = "ENABLED";
    FD1P3AX array_255___i1102 (.D(array_0__7__N_3001[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[118] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1102.GSR = "ENABLED";
    FD1P3AX array_255___i1103 (.D(array_0__7__N_3001[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[118] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1103.GSR = "ENABLED";
    FD1P3AX array_255___i1104 (.D(array_0__7__N_3001[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[118] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1104.GSR = "ENABLED";
    FD1P3AX array_255___i1105 (.D(array_0__7__N_2993[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[117] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1105.GSR = "ENABLED";
    FD1P3AX array_255___i1106 (.D(array_0__7__N_2993[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[117] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1106.GSR = "ENABLED";
    FD1P3AX array_255___i1107 (.D(array_0__7__N_2993[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[117] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1107.GSR = "ENABLED";
    FD1P3AX array_255___i1108 (.D(array_0__7__N_2993[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[117] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1108.GSR = "ENABLED";
    FD1P3AX array_255___i1109 (.D(array_0__7__N_2993[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[117] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1109.GSR = "ENABLED";
    FD1P3AX array_255___i1110 (.D(array_0__7__N_2993[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[117] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1110.GSR = "ENABLED";
    FD1P3AX array_255___i1111 (.D(array_0__7__N_2993[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[117] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1111.GSR = "ENABLED";
    FD1P3AX array_255___i1112 (.D(array_0__7__N_2993[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[117] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1112.GSR = "ENABLED";
    FD1P3AX array_255___i1113 (.D(array_0__7__N_2985[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[116] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1113.GSR = "ENABLED";
    FD1P3AX array_255___i1114 (.D(array_0__7__N_2985[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[116] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1114.GSR = "ENABLED";
    FD1P3AX array_255___i1115 (.D(array_0__7__N_2985[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[116] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1115.GSR = "ENABLED";
    FD1P3AX array_255___i1116 (.D(array_0__7__N_2985[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[116] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1116.GSR = "ENABLED";
    FD1P3AX array_255___i1117 (.D(array_0__7__N_2985[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[116] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1117.GSR = "ENABLED";
    FD1P3AX array_255___i1118 (.D(array_0__7__N_2985[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[116] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1118.GSR = "ENABLED";
    FD1P3AX array_255___i1119 (.D(array_0__7__N_2985[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[116] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1119.GSR = "ENABLED";
    FD1P3AX array_255___i1120 (.D(array_0__7__N_2985[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[116] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1120.GSR = "ENABLED";
    FD1P3AX array_255___i1121 (.D(array_0__7__N_2977[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[115] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1121.GSR = "ENABLED";
    FD1P3AX array_255___i1122 (.D(array_0__7__N_2977[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[115] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1122.GSR = "ENABLED";
    FD1P3AX array_255___i1123 (.D(array_0__7__N_2977[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[115] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1123.GSR = "ENABLED";
    FD1P3AX array_255___i1124 (.D(array_0__7__N_2977[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[115] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1124.GSR = "ENABLED";
    FD1P3AX array_255___i1125 (.D(array_0__7__N_2977[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[115] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1125.GSR = "ENABLED";
    FD1P3AX array_255___i1126 (.D(array_0__7__N_2977[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[115] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1126.GSR = "ENABLED";
    FD1P3AX array_255___i1127 (.D(array_0__7__N_2977[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[115] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1127.GSR = "ENABLED";
    FD1P3AX array_255___i1128 (.D(array_0__7__N_2977[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[115] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1128.GSR = "ENABLED";
    FD1P3AX array_255___i1129 (.D(array_0__7__N_2969[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[114] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1129.GSR = "ENABLED";
    FD1P3AX array_255___i1130 (.D(array_0__7__N_2969[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[114] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1130.GSR = "ENABLED";
    FD1P3AX array_255___i1131 (.D(array_0__7__N_2969[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[114] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1131.GSR = "ENABLED";
    FD1P3AX array_255___i1132 (.D(array_0__7__N_2969[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[114] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1132.GSR = "ENABLED";
    FD1P3AX array_255___i1133 (.D(array_0__7__N_2969[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[114] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1133.GSR = "ENABLED";
    FD1P3AX array_255___i1134 (.D(array_0__7__N_2969[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[114] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1134.GSR = "ENABLED";
    FD1P3AX array_255___i1135 (.D(array_0__7__N_2969[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[114] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1135.GSR = "ENABLED";
    FD1P3AX array_255___i1136 (.D(array_0__7__N_2969[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[114] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1136.GSR = "ENABLED";
    FD1P3AX array_255___i1137 (.D(array_0__7__N_2961[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[113] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1137.GSR = "ENABLED";
    FD1P3AX array_255___i1138 (.D(array_0__7__N_2961[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[113] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1138.GSR = "ENABLED";
    FD1P3AX array_255___i1139 (.D(array_0__7__N_2961[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[113] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1139.GSR = "ENABLED";
    FD1P3AX array_255___i1140 (.D(array_0__7__N_2961[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[113] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1140.GSR = "ENABLED";
    FD1P3AX array_255___i1141 (.D(array_0__7__N_2961[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[113] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1141.GSR = "ENABLED";
    FD1P3AX array_255___i1142 (.D(array_0__7__N_2961[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[113] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1142.GSR = "ENABLED";
    FD1P3AX array_255___i1143 (.D(array_0__7__N_2961[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[113] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1143.GSR = "ENABLED";
    FD1P3AX array_255___i1144 (.D(array_0__7__N_2961[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[113] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1144.GSR = "ENABLED";
    FD1P3AX array_255___i1145 (.D(array_0__7__N_2953[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[112] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1145.GSR = "ENABLED";
    FD1P3AX array_255___i1146 (.D(array_0__7__N_2953[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[112] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1146.GSR = "ENABLED";
    FD1P3AX array_255___i1147 (.D(array_0__7__N_2953[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[112] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1147.GSR = "ENABLED";
    FD1P3AX array_255___i1148 (.D(array_0__7__N_2953[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[112] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1148.GSR = "ENABLED";
    FD1P3AX array_255___i1149 (.D(array_0__7__N_2953[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[112] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1149.GSR = "ENABLED";
    FD1P3AX array_255___i1150 (.D(array_0__7__N_2953[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[112] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1150.GSR = "ENABLED";
    FD1P3AX array_255___i1151 (.D(array_0__7__N_2953[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[112] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1151.GSR = "ENABLED";
    FD1P3AX array_255___i1152 (.D(array_0__7__N_2953[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[112] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1152.GSR = "ENABLED";
    FD1P3AX array_255___i1153 (.D(array_0__7__N_2945[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[111] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1153.GSR = "ENABLED";
    FD1P3AX array_255___i1154 (.D(array_0__7__N_2945[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[111] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1154.GSR = "ENABLED";
    FD1P3AX array_255___i1155 (.D(array_0__7__N_2945[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[111] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1155.GSR = "ENABLED";
    FD1P3AX array_255___i1156 (.D(array_0__7__N_2945[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[111] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1156.GSR = "ENABLED";
    FD1P3AX array_255___i1157 (.D(array_0__7__N_2945[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[111] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1157.GSR = "ENABLED";
    FD1P3AX array_255___i1158 (.D(array_0__7__N_2945[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[111] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1158.GSR = "ENABLED";
    FD1P3AX array_255___i1159 (.D(array_0__7__N_2945[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[111] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1159.GSR = "ENABLED";
    FD1P3AX array_255___i1160 (.D(array_0__7__N_2945[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[111] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1160.GSR = "ENABLED";
    FD1P3AX array_255___i1161 (.D(array_0__7__N_2937[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[110] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1161.GSR = "ENABLED";
    FD1P3AX array_255___i1162 (.D(array_0__7__N_2937[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[110] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1162.GSR = "ENABLED";
    FD1P3AX array_255___i1163 (.D(array_0__7__N_2937[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[110] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1163.GSR = "ENABLED";
    FD1P3AX array_255___i1164 (.D(array_0__7__N_2937[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[110] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1164.GSR = "ENABLED";
    FD1P3AX array_255___i1165 (.D(array_0__7__N_2937[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[110] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1165.GSR = "ENABLED";
    FD1P3AX array_255___i1166 (.D(array_0__7__N_2937[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[110] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1166.GSR = "ENABLED";
    FD1P3AX array_255___i1167 (.D(array_0__7__N_2937[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[110] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1167.GSR = "ENABLED";
    FD1P3AX array_255___i1168 (.D(array_0__7__N_2937[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[110] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1168.GSR = "ENABLED";
    FD1P3AX array_255___i1169 (.D(array_0__7__N_2929[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[109] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1169.GSR = "ENABLED";
    FD1P3AX array_255___i1170 (.D(array_0__7__N_2929[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[109] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1170.GSR = "ENABLED";
    FD1P3AX array_255___i1171 (.D(array_0__7__N_2929[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[109] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1171.GSR = "ENABLED";
    FD1P3AX array_255___i1172 (.D(array_0__7__N_2929[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[109] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1172.GSR = "ENABLED";
    FD1P3AX array_255___i1173 (.D(array_0__7__N_2929[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[109] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1173.GSR = "ENABLED";
    FD1P3AX array_255___i1174 (.D(array_0__7__N_2929[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[109] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1174.GSR = "ENABLED";
    FD1P3AX array_255___i1175 (.D(array_0__7__N_2929[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[109] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1175.GSR = "ENABLED";
    FD1P3AX array_255___i1176 (.D(array_0__7__N_2929[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[109] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1176.GSR = "ENABLED";
    FD1P3AX array_255___i1177 (.D(array_0__7__N_2921[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[108] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1177.GSR = "ENABLED";
    FD1P3AX array_255___i1178 (.D(array_0__7__N_2921[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[108] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1178.GSR = "ENABLED";
    FD1P3AX array_255___i1179 (.D(array_0__7__N_2921[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[108] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1179.GSR = "ENABLED";
    FD1P3AX array_255___i1180 (.D(array_0__7__N_2921[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[108] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1180.GSR = "ENABLED";
    FD1P3AX array_255___i1181 (.D(array_0__7__N_2921[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[108] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1181.GSR = "ENABLED";
    FD1P3AX array_255___i1182 (.D(array_0__7__N_2921[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[108] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1182.GSR = "ENABLED";
    FD1P3AX array_255___i1183 (.D(array_0__7__N_2921[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[108] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1183.GSR = "ENABLED";
    FD1P3AX array_255___i1184 (.D(array_0__7__N_2921[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[108] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1184.GSR = "ENABLED";
    FD1P3AX array_255___i1185 (.D(array_0__7__N_2913[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[107] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1185.GSR = "ENABLED";
    FD1P3AX array_255___i1186 (.D(array_0__7__N_2913[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[107] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1186.GSR = "ENABLED";
    FD1P3AX array_255___i1187 (.D(array_0__7__N_2913[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[107] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1187.GSR = "ENABLED";
    FD1P3AX array_255___i1188 (.D(array_0__7__N_2913[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[107] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1188.GSR = "ENABLED";
    FD1P3AX array_255___i1189 (.D(array_0__7__N_2913[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[107] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1189.GSR = "ENABLED";
    FD1P3AX array_255___i1190 (.D(array_0__7__N_2913[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[107] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1190.GSR = "ENABLED";
    FD1P3AX array_255___i1191 (.D(array_0__7__N_2913[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[107] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1191.GSR = "ENABLED";
    FD1P3AX array_255___i1192 (.D(array_0__7__N_2913[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[107] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1192.GSR = "ENABLED";
    FD1P3AX array_255___i1193 (.D(array_0__7__N_2905[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[106] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1193.GSR = "ENABLED";
    FD1P3AX array_255___i1194 (.D(array_0__7__N_2905[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[106] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1194.GSR = "ENABLED";
    FD1P3AX array_255___i1195 (.D(array_0__7__N_2905[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[106] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1195.GSR = "ENABLED";
    FD1P3AX array_255___i1196 (.D(array_0__7__N_2905[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[106] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1196.GSR = "ENABLED";
    FD1P3AX array_255___i1197 (.D(array_0__7__N_2905[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[106] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1197.GSR = "ENABLED";
    FD1P3AX array_255___i1198 (.D(array_0__7__N_2905[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[106] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1198.GSR = "ENABLED";
    FD1P3AX array_255___i1199 (.D(array_0__7__N_2905[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[106] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1199.GSR = "ENABLED";
    FD1P3AX array_255___i1200 (.D(array_0__7__N_2905[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[106] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1200.GSR = "ENABLED";
    FD1P3AX array_255___i1201 (.D(array_0__7__N_2897[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[105] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1201.GSR = "ENABLED";
    FD1P3AX array_255___i1202 (.D(array_0__7__N_2897[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[105] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1202.GSR = "ENABLED";
    FD1P3AX array_255___i1203 (.D(array_0__7__N_2897[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[105] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1203.GSR = "ENABLED";
    FD1P3AX array_255___i1204 (.D(array_0__7__N_2897[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[105] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1204.GSR = "ENABLED";
    FD1P3AX array_255___i1205 (.D(array_0__7__N_2897[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[105] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1205.GSR = "ENABLED";
    FD1P3AX array_255___i1206 (.D(array_0__7__N_2897[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[105] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1206.GSR = "ENABLED";
    FD1P3AX array_255___i1207 (.D(array_0__7__N_2897[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[105] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1207.GSR = "ENABLED";
    FD1P3AX array_255___i1208 (.D(array_0__7__N_2897[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[105] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1208.GSR = "ENABLED";
    FD1P3AX array_255___i1209 (.D(array_0__7__N_2889[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[104] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1209.GSR = "ENABLED";
    FD1P3AX array_255___i1210 (.D(array_0__7__N_2889[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[104] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1210.GSR = "ENABLED";
    FD1P3AX array_255___i1211 (.D(array_0__7__N_2889[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[104] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1211.GSR = "ENABLED";
    FD1P3AX array_255___i1212 (.D(array_0__7__N_2889[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[104] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1212.GSR = "ENABLED";
    FD1P3AX array_255___i1213 (.D(array_0__7__N_2889[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[104] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1213.GSR = "ENABLED";
    FD1P3AX array_255___i1214 (.D(array_0__7__N_2889[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[104] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1214.GSR = "ENABLED";
    FD1P3AX array_255___i1215 (.D(array_0__7__N_2889[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[104] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1215.GSR = "ENABLED";
    FD1P3AX array_255___i1216 (.D(array_0__7__N_2889[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[104] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1216.GSR = "ENABLED";
    FD1P3AX array_255___i1217 (.D(array_0__7__N_2881[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[103] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1217.GSR = "ENABLED";
    FD1P3AX array_255___i1218 (.D(array_0__7__N_2881[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[103] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1218.GSR = "ENABLED";
    FD1P3AX array_255___i1219 (.D(array_0__7__N_2881[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[103] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1219.GSR = "ENABLED";
    FD1P3AX array_255___i1220 (.D(array_0__7__N_2881[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[103] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1220.GSR = "ENABLED";
    FD1P3AX array_255___i1221 (.D(array_0__7__N_2881[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[103] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1221.GSR = "ENABLED";
    FD1P3AX array_255___i1222 (.D(array_0__7__N_2881[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[103] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1222.GSR = "ENABLED";
    FD1P3AX array_255___i1223 (.D(array_0__7__N_2881[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[103] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1223.GSR = "ENABLED";
    FD1P3AX array_255___i1224 (.D(array_0__7__N_2881[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[103] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1224.GSR = "ENABLED";
    FD1P3AX array_255___i1225 (.D(array_0__7__N_2873[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[102] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1225.GSR = "ENABLED";
    FD1P3AX array_255___i1226 (.D(array_0__7__N_2873[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[102] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1226.GSR = "ENABLED";
    FD1P3AX array_255___i1227 (.D(array_0__7__N_2873[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[102] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1227.GSR = "ENABLED";
    FD1P3AX array_255___i1228 (.D(array_0__7__N_2873[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[102] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1228.GSR = "ENABLED";
    FD1P3AX array_255___i1229 (.D(array_0__7__N_2873[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[102] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1229.GSR = "ENABLED";
    FD1P3AX array_255___i1230 (.D(array_0__7__N_2873[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[102] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1230.GSR = "ENABLED";
    FD1P3AX array_255___i1231 (.D(array_0__7__N_2873[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[102] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1231.GSR = "ENABLED";
    FD1P3AX array_255___i1232 (.D(array_0__7__N_2873[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[102] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1232.GSR = "ENABLED";
    FD1P3AX array_255___i1233 (.D(array_0__7__N_2865[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[101] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1233.GSR = "ENABLED";
    FD1P3AX array_255___i1234 (.D(array_0__7__N_2865[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[101] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1234.GSR = "ENABLED";
    FD1P3AX array_255___i1235 (.D(array_0__7__N_2865[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[101] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1235.GSR = "ENABLED";
    FD1P3AX array_255___i1236 (.D(array_0__7__N_2865[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[101] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1236.GSR = "ENABLED";
    FD1P3AX array_255___i1237 (.D(array_0__7__N_2865[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[101] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1237.GSR = "ENABLED";
    FD1P3AX array_255___i1238 (.D(array_0__7__N_2865[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[101] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1238.GSR = "ENABLED";
    FD1P3AX array_255___i1239 (.D(array_0__7__N_2865[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[101] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1239.GSR = "ENABLED";
    FD1P3AX array_255___i1240 (.D(array_0__7__N_2865[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[101] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1240.GSR = "ENABLED";
    FD1P3AX array_255___i1241 (.D(array_0__7__N_2857[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[100] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1241.GSR = "ENABLED";
    FD1P3AX array_255___i1242 (.D(array_0__7__N_2857[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[100] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1242.GSR = "ENABLED";
    FD1P3AX array_255___i1243 (.D(array_0__7__N_2857[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[100] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1243.GSR = "ENABLED";
    FD1P3AX array_255___i1244 (.D(array_0__7__N_2857[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[100] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1244.GSR = "ENABLED";
    FD1P3AX array_255___i1245 (.D(array_0__7__N_2857[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[100] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1245.GSR = "ENABLED";
    FD1P3AX array_255___i1246 (.D(array_0__7__N_2857[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[100] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1246.GSR = "ENABLED";
    FD1P3AX array_255___i1247 (.D(array_0__7__N_2857[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[100] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1247.GSR = "ENABLED";
    FD1P3AX array_255___i1248 (.D(array_0__7__N_2857[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[100] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1248.GSR = "ENABLED";
    FD1P3AX array_255___i1249 (.D(array_0__7__N_2849[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[99] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1249.GSR = "ENABLED";
    FD1P3AX array_255___i1250 (.D(array_0__7__N_2849[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[99] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1250.GSR = "ENABLED";
    FD1P3AX array_255___i1251 (.D(array_0__7__N_2849[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[99] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1251.GSR = "ENABLED";
    FD1P3AX array_255___i1252 (.D(array_0__7__N_2849[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[99] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1252.GSR = "ENABLED";
    FD1P3AX array_255___i1253 (.D(array_0__7__N_2849[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[99] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1253.GSR = "ENABLED";
    FD1P3AX array_255___i1254 (.D(array_0__7__N_2849[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[99] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1254.GSR = "ENABLED";
    FD1P3AX array_255___i1255 (.D(array_0__7__N_2849[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[99] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1255.GSR = "ENABLED";
    FD1P3AX array_255___i1256 (.D(array_0__7__N_2849[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[99] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1256.GSR = "ENABLED";
    FD1P3AX array_255___i1257 (.D(array_0__7__N_2841[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[98] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1257.GSR = "ENABLED";
    FD1P3AX array_255___i1258 (.D(array_0__7__N_2841[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[98] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1258.GSR = "ENABLED";
    FD1P3AX array_255___i1259 (.D(array_0__7__N_2841[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[98] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1259.GSR = "ENABLED";
    FD1P3AX array_255___i1260 (.D(array_0__7__N_2841[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[98] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1260.GSR = "ENABLED";
    FD1P3AX array_255___i1261 (.D(array_0__7__N_2841[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[98] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1261.GSR = "ENABLED";
    FD1P3AX array_255___i1262 (.D(array_0__7__N_2841[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[98] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1262.GSR = "ENABLED";
    FD1P3AX array_255___i1263 (.D(array_0__7__N_2841[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[98] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1263.GSR = "ENABLED";
    FD1P3AX array_255___i1264 (.D(array_0__7__N_2841[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[98] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1264.GSR = "ENABLED";
    FD1P3AX array_255___i1265 (.D(array_0__7__N_2833[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[97] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1265.GSR = "ENABLED";
    FD1P3AX array_255___i1266 (.D(array_0__7__N_2833[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[97] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1266.GSR = "ENABLED";
    FD1P3AX array_255___i1267 (.D(array_0__7__N_2833[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[97] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1267.GSR = "ENABLED";
    FD1P3AX array_255___i1268 (.D(array_0__7__N_2833[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[97] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1268.GSR = "ENABLED";
    FD1P3AX array_255___i1269 (.D(array_0__7__N_2833[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[97] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1269.GSR = "ENABLED";
    FD1P3AX array_255___i1270 (.D(array_0__7__N_2833[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[97] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1270.GSR = "ENABLED";
    FD1P3AX array_255___i1271 (.D(array_0__7__N_2833[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[97] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1271.GSR = "ENABLED";
    FD1P3AX array_255___i1272 (.D(array_0__7__N_2833[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[97] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1272.GSR = "ENABLED";
    FD1P3AX array_255___i1273 (.D(array_0__7__N_2825[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[96] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1273.GSR = "ENABLED";
    FD1P3AX array_255___i1274 (.D(array_0__7__N_2825[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[96] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1274.GSR = "ENABLED";
    FD1P3AX array_255___i1275 (.D(array_0__7__N_2825[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[96] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1275.GSR = "ENABLED";
    FD1P3AX array_255___i1276 (.D(array_0__7__N_2825[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[96] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1276.GSR = "ENABLED";
    FD1P3AX array_255___i1277 (.D(array_0__7__N_2825[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[96] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1277.GSR = "ENABLED";
    FD1P3AX array_255___i1278 (.D(array_0__7__N_2825[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[96] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1278.GSR = "ENABLED";
    FD1P3AX array_255___i1279 (.D(array_0__7__N_2825[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[96] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1279.GSR = "ENABLED";
    FD1P3AX array_255___i1280 (.D(array_0__7__N_2825[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[96] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1280.GSR = "ENABLED";
    FD1P3AX array_255___i1281 (.D(array_0__7__N_2817[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[95] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1281.GSR = "ENABLED";
    FD1P3AX array_255___i1282 (.D(array_0__7__N_2817[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[95] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1282.GSR = "ENABLED";
    FD1P3AX array_255___i1283 (.D(array_0__7__N_2817[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[95] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1283.GSR = "ENABLED";
    FD1P3AX array_255___i1284 (.D(array_0__7__N_2817[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[95] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1284.GSR = "ENABLED";
    FD1P3AX array_255___i1285 (.D(array_0__7__N_2817[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[95] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1285.GSR = "ENABLED";
    FD1P3AX array_255___i1286 (.D(array_0__7__N_2817[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[95] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1286.GSR = "ENABLED";
    FD1P3AX array_255___i1287 (.D(array_0__7__N_2817[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[95] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1287.GSR = "ENABLED";
    FD1P3AX array_255___i1288 (.D(array_0__7__N_2817[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[95] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1288.GSR = "ENABLED";
    FD1P3AX array_255___i1289 (.D(array_0__7__N_2809[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[94] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1289.GSR = "ENABLED";
    FD1P3AX array_255___i1290 (.D(array_0__7__N_2809[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[94] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1290.GSR = "ENABLED";
    FD1P3AX array_255___i1291 (.D(array_0__7__N_2809[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[94] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1291.GSR = "ENABLED";
    FD1P3AX array_255___i1292 (.D(array_0__7__N_2809[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[94] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1292.GSR = "ENABLED";
    FD1P3AX array_255___i1293 (.D(array_0__7__N_2809[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[94] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1293.GSR = "ENABLED";
    FD1P3AX array_255___i1294 (.D(array_0__7__N_2809[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[94] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1294.GSR = "ENABLED";
    FD1P3AX array_255___i1295 (.D(array_0__7__N_2809[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[94] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1295.GSR = "ENABLED";
    FD1P3AX array_255___i1296 (.D(array_0__7__N_2809[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[94] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1296.GSR = "ENABLED";
    FD1P3AX array_255___i1297 (.D(array_0__7__N_2801[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[93] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1297.GSR = "ENABLED";
    FD1P3AX array_255___i1298 (.D(array_0__7__N_2801[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[93] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1298.GSR = "ENABLED";
    FD1P3AX array_255___i1299 (.D(array_0__7__N_2801[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[93] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1299.GSR = "ENABLED";
    FD1P3AX array_255___i1300 (.D(array_0__7__N_2801[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[93] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1300.GSR = "ENABLED";
    FD1P3AX array_255___i1301 (.D(array_0__7__N_2801[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[93] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1301.GSR = "ENABLED";
    FD1P3AX array_255___i1302 (.D(array_0__7__N_2801[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[93] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1302.GSR = "ENABLED";
    FD1P3AX array_255___i1303 (.D(array_0__7__N_2801[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[93] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1303.GSR = "ENABLED";
    FD1P3AX array_255___i1304 (.D(array_0__7__N_2801[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[93] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1304.GSR = "ENABLED";
    FD1P3AX array_255___i1305 (.D(array_0__7__N_2793[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[92] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1305.GSR = "ENABLED";
    FD1P3AX array_255___i1306 (.D(array_0__7__N_2793[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[92] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1306.GSR = "ENABLED";
    FD1P3AX array_255___i1307 (.D(array_0__7__N_2793[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[92] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1307.GSR = "ENABLED";
    FD1P3AX array_255___i1308 (.D(array_0__7__N_2793[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[92] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1308.GSR = "ENABLED";
    FD1P3AX array_255___i1309 (.D(array_0__7__N_2793[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[92] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1309.GSR = "ENABLED";
    FD1P3AX array_255___i1310 (.D(array_0__7__N_2793[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[92] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1310.GSR = "ENABLED";
    FD1P3AX array_255___i1311 (.D(array_0__7__N_2793[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[92] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1311.GSR = "ENABLED";
    FD1P3AX array_255___i1312 (.D(array_0__7__N_2793[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[92] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1312.GSR = "ENABLED";
    FD1P3AX array_255___i1313 (.D(array_0__7__N_2785[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[91] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1313.GSR = "ENABLED";
    FD1P3AX array_255___i1314 (.D(array_0__7__N_2785[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[91] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1314.GSR = "ENABLED";
    FD1P3AX array_255___i1315 (.D(array_0__7__N_2785[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[91] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1315.GSR = "ENABLED";
    FD1P3AX array_255___i1316 (.D(array_0__7__N_2785[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[91] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1316.GSR = "ENABLED";
    FD1P3AX array_255___i1317 (.D(array_0__7__N_2785[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[91] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1317.GSR = "ENABLED";
    FD1P3AX array_255___i1318 (.D(array_0__7__N_2785[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[91] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1318.GSR = "ENABLED";
    FD1P3AX array_255___i1319 (.D(array_0__7__N_2785[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[91] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1319.GSR = "ENABLED";
    FD1P3AX array_255___i1320 (.D(array_0__7__N_2785[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[91] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1320.GSR = "ENABLED";
    FD1P3AX array_255___i1321 (.D(array_0__7__N_2777[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[90] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1321.GSR = "ENABLED";
    FD1P3AX array_255___i1322 (.D(array_0__7__N_2777[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[90] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1322.GSR = "ENABLED";
    FD1P3AX array_255___i1323 (.D(array_0__7__N_2777[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[90] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1323.GSR = "ENABLED";
    FD1P3AX array_255___i1324 (.D(array_0__7__N_2777[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[90] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1324.GSR = "ENABLED";
    FD1P3AX array_255___i1325 (.D(array_0__7__N_2777[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[90] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1325.GSR = "ENABLED";
    FD1P3AX array_255___i1326 (.D(array_0__7__N_2777[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[90] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1326.GSR = "ENABLED";
    FD1P3AX array_255___i1327 (.D(array_0__7__N_2777[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[90] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1327.GSR = "ENABLED";
    FD1P3AX array_255___i1328 (.D(array_0__7__N_2777[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[90] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1328.GSR = "ENABLED";
    FD1P3AX array_255___i1329 (.D(array_0__7__N_2769[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[89] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1329.GSR = "ENABLED";
    FD1P3AX array_255___i1330 (.D(array_0__7__N_2769[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[89] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1330.GSR = "ENABLED";
    FD1P3AX array_255___i1331 (.D(array_0__7__N_2769[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[89] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1331.GSR = "ENABLED";
    FD1P3AX array_255___i1332 (.D(array_0__7__N_2769[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[89] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1332.GSR = "ENABLED";
    FD1P3AX array_255___i1333 (.D(array_0__7__N_2769[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[89] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1333.GSR = "ENABLED";
    FD1P3AX array_255___i1334 (.D(array_0__7__N_2769[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[89] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1334.GSR = "ENABLED";
    FD1P3AX array_255___i1335 (.D(array_0__7__N_2769[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[89] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1335.GSR = "ENABLED";
    FD1P3AX array_255___i1336 (.D(array_0__7__N_2769[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[89] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1336.GSR = "ENABLED";
    FD1P3AX array_255___i1337 (.D(array_0__7__N_2761[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[88] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1337.GSR = "ENABLED";
    FD1P3AX array_255___i1338 (.D(array_0__7__N_2761[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[88] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1338.GSR = "ENABLED";
    FD1P3AX array_255___i1339 (.D(array_0__7__N_2761[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[88] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1339.GSR = "ENABLED";
    FD1P3AX array_255___i1340 (.D(array_0__7__N_2761[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[88] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1340.GSR = "ENABLED";
    FD1P3AX array_255___i1341 (.D(array_0__7__N_2761[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[88] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1341.GSR = "ENABLED";
    FD1P3AX array_255___i1342 (.D(array_0__7__N_2761[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[88] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1342.GSR = "ENABLED";
    FD1P3AX array_255___i1343 (.D(array_0__7__N_2761[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[88] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1343.GSR = "ENABLED";
    FD1P3AX array_255___i1344 (.D(array_0__7__N_2761[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[88] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1344.GSR = "ENABLED";
    FD1P3AX array_255___i1345 (.D(array_0__7__N_2753[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[87] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1345.GSR = "ENABLED";
    FD1P3AX array_255___i1346 (.D(array_0__7__N_2753[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[87] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1346.GSR = "ENABLED";
    FD1P3AX array_255___i1347 (.D(array_0__7__N_2753[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[87] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1347.GSR = "ENABLED";
    FD1P3AX array_255___i1348 (.D(array_0__7__N_2753[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[87] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1348.GSR = "ENABLED";
    FD1P3AX array_255___i1349 (.D(array_0__7__N_2753[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[87] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1349.GSR = "ENABLED";
    FD1P3AX array_255___i1350 (.D(array_0__7__N_2753[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[87] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1350.GSR = "ENABLED";
    FD1P3AX array_255___i1351 (.D(array_0__7__N_2753[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[87] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1351.GSR = "ENABLED";
    FD1P3AX array_255___i1352 (.D(array_0__7__N_2753[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[87] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1352.GSR = "ENABLED";
    FD1P3AX array_255___i1353 (.D(array_0__7__N_2745[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[86] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1353.GSR = "ENABLED";
    FD1P3AX array_255___i1354 (.D(array_0__7__N_2745[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[86] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1354.GSR = "ENABLED";
    FD1P3AX array_255___i1355 (.D(array_0__7__N_2745[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[86] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1355.GSR = "ENABLED";
    FD1P3AX array_255___i1356 (.D(array_0__7__N_2745[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[86] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1356.GSR = "ENABLED";
    FD1P3AX array_255___i1357 (.D(array_0__7__N_2745[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[86] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1357.GSR = "ENABLED";
    FD1P3AX array_255___i1358 (.D(array_0__7__N_2745[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[86] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1358.GSR = "ENABLED";
    FD1P3AX array_255___i1359 (.D(array_0__7__N_2745[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[86] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1359.GSR = "ENABLED";
    FD1P3AX array_255___i1360 (.D(array_0__7__N_2745[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[86] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1360.GSR = "ENABLED";
    FD1P3AX array_255___i1361 (.D(array_0__7__N_2737[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[85] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1361.GSR = "ENABLED";
    FD1P3AX array_255___i1362 (.D(array_0__7__N_2737[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[85] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1362.GSR = "ENABLED";
    FD1P3AX array_255___i1363 (.D(array_0__7__N_2737[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[85] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1363.GSR = "ENABLED";
    FD1P3AX array_255___i1364 (.D(array_0__7__N_2737[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[85] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1364.GSR = "ENABLED";
    FD1P3AX array_255___i1365 (.D(array_0__7__N_2737[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[85] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1365.GSR = "ENABLED";
    FD1P3AX array_255___i1366 (.D(array_0__7__N_2737[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[85] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1366.GSR = "ENABLED";
    FD1P3AX array_255___i1367 (.D(array_0__7__N_2737[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[85] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1367.GSR = "ENABLED";
    FD1P3AX array_255___i1368 (.D(array_0__7__N_2737[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[85] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1368.GSR = "ENABLED";
    FD1P3AX array_255___i1369 (.D(array_0__7__N_2729[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[84] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1369.GSR = "ENABLED";
    FD1P3AX array_255___i1370 (.D(array_0__7__N_2729[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[84] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1370.GSR = "ENABLED";
    FD1P3AX array_255___i1371 (.D(array_0__7__N_2729[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[84] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1371.GSR = "ENABLED";
    FD1P3AX array_255___i1372 (.D(array_0__7__N_2729[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[84] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1372.GSR = "ENABLED";
    FD1P3AX array_255___i1373 (.D(array_0__7__N_2729[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[84] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1373.GSR = "ENABLED";
    FD1P3AX array_255___i1374 (.D(array_0__7__N_2729[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[84] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1374.GSR = "ENABLED";
    FD1P3AX array_255___i1375 (.D(array_0__7__N_2729[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[84] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1375.GSR = "ENABLED";
    FD1P3AX array_255___i1376 (.D(array_0__7__N_2729[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[84] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1376.GSR = "ENABLED";
    FD1P3AX array_255___i1377 (.D(array_0__7__N_2721[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[83] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1377.GSR = "ENABLED";
    FD1P3AX array_255___i1378 (.D(array_0__7__N_2721[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[83] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1378.GSR = "ENABLED";
    FD1P3AX array_255___i1379 (.D(array_0__7__N_2721[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[83] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1379.GSR = "ENABLED";
    FD1P3AX array_255___i1380 (.D(array_0__7__N_2721[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[83] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1380.GSR = "ENABLED";
    FD1P3AX array_255___i1381 (.D(array_0__7__N_2721[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[83] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1381.GSR = "ENABLED";
    FD1P3AX array_255___i1382 (.D(array_0__7__N_2721[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[83] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1382.GSR = "ENABLED";
    FD1P3AX array_255___i1383 (.D(array_0__7__N_2721[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[83] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1383.GSR = "ENABLED";
    FD1P3AX array_255___i1384 (.D(array_0__7__N_2721[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[83] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1384.GSR = "ENABLED";
    FD1P3AX array_255___i1385 (.D(array_0__7__N_2713[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[82] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1385.GSR = "ENABLED";
    FD1P3AX array_255___i1386 (.D(array_0__7__N_2713[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[82] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1386.GSR = "ENABLED";
    FD1P3AX array_255___i1387 (.D(array_0__7__N_2713[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[82] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1387.GSR = "ENABLED";
    FD1P3AX array_255___i1388 (.D(array_0__7__N_2713[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[82] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1388.GSR = "ENABLED";
    FD1P3AX array_255___i1389 (.D(array_0__7__N_2713[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[82] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1389.GSR = "ENABLED";
    FD1P3AX array_255___i1390 (.D(array_0__7__N_2713[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[82] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1390.GSR = "ENABLED";
    FD1P3AX array_255___i1391 (.D(array_0__7__N_2713[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[82] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1391.GSR = "ENABLED";
    FD1P3AX array_255___i1392 (.D(array_0__7__N_2713[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[82] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1392.GSR = "ENABLED";
    FD1P3AX array_255___i1393 (.D(array_0__7__N_2705[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[81] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1393.GSR = "ENABLED";
    FD1P3AX array_255___i1394 (.D(array_0__7__N_2705[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[81] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1394.GSR = "ENABLED";
    FD1P3AX array_255___i1395 (.D(array_0__7__N_2705[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[81] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1395.GSR = "ENABLED";
    FD1P3AX array_255___i1396 (.D(array_0__7__N_2705[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[81] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1396.GSR = "ENABLED";
    FD1P3AX array_255___i1397 (.D(array_0__7__N_2705[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[81] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1397.GSR = "ENABLED";
    FD1P3AX array_255___i1398 (.D(array_0__7__N_2705[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[81] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1398.GSR = "ENABLED";
    FD1P3AX array_255___i1399 (.D(array_0__7__N_2705[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[81] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1399.GSR = "ENABLED";
    FD1P3AX array_255___i1400 (.D(array_0__7__N_2705[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[81] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1400.GSR = "ENABLED";
    FD1P3AX array_255___i1401 (.D(array_0__7__N_2697[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[80] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1401.GSR = "ENABLED";
    FD1P3AX array_255___i1402 (.D(array_0__7__N_2697[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[80] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1402.GSR = "ENABLED";
    FD1P3AX array_255___i1403 (.D(array_0__7__N_2697[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[80] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1403.GSR = "ENABLED";
    FD1P3AX array_255___i1404 (.D(array_0__7__N_2697[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[80] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1404.GSR = "ENABLED";
    FD1P3AX array_255___i1405 (.D(array_0__7__N_2697[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[80] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1405.GSR = "ENABLED";
    FD1P3AX array_255___i1406 (.D(array_0__7__N_2697[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[80] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1406.GSR = "ENABLED";
    FD1P3AX array_255___i1407 (.D(array_0__7__N_2697[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[80] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1407.GSR = "ENABLED";
    FD1P3AX array_255___i1408 (.D(array_0__7__N_2697[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[80] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1408.GSR = "ENABLED";
    FD1P3AX array_255___i1409 (.D(array_0__7__N_2689[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[79] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1409.GSR = "ENABLED";
    FD1P3AX array_255___i1410 (.D(array_0__7__N_2689[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[79] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1410.GSR = "ENABLED";
    FD1P3AX array_255___i1411 (.D(array_0__7__N_2689[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[79] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1411.GSR = "ENABLED";
    FD1P3AX array_255___i1412 (.D(array_0__7__N_2689[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[79] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1412.GSR = "ENABLED";
    FD1P3AX array_255___i1413 (.D(array_0__7__N_2689[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[79] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1413.GSR = "ENABLED";
    FD1P3AX array_255___i1414 (.D(array_0__7__N_2689[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[79] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1414.GSR = "ENABLED";
    FD1P3AX array_255___i1415 (.D(array_0__7__N_2689[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[79] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1415.GSR = "ENABLED";
    FD1P3AX array_255___i1416 (.D(array_0__7__N_2689[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[79] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1416.GSR = "ENABLED";
    FD1P3AX array_255___i1417 (.D(array_0__7__N_2681[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[78] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1417.GSR = "ENABLED";
    FD1P3AX array_255___i1418 (.D(array_0__7__N_2681[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[78] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1418.GSR = "ENABLED";
    FD1P3AX array_255___i1419 (.D(array_0__7__N_2681[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[78] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1419.GSR = "ENABLED";
    FD1P3AX array_255___i1420 (.D(array_0__7__N_2681[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[78] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1420.GSR = "ENABLED";
    FD1P3AX array_255___i1421 (.D(array_0__7__N_2681[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[78] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1421.GSR = "ENABLED";
    FD1P3AX array_255___i1422 (.D(array_0__7__N_2681[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[78] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1422.GSR = "ENABLED";
    FD1P3AX array_255___i1423 (.D(array_0__7__N_2681[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[78] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1423.GSR = "ENABLED";
    FD1P3AX array_255___i1424 (.D(array_0__7__N_2681[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[78] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1424.GSR = "ENABLED";
    FD1P3AX array_255___i1425 (.D(array_0__7__N_2673[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[77] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1425.GSR = "ENABLED";
    FD1P3AX array_255___i1426 (.D(array_0__7__N_2673[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[77] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1426.GSR = "ENABLED";
    FD1P3AX array_255___i1427 (.D(array_0__7__N_2673[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[77] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1427.GSR = "ENABLED";
    FD1P3AX array_255___i1428 (.D(array_0__7__N_2673[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[77] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1428.GSR = "ENABLED";
    FD1P3AX array_255___i1429 (.D(array_0__7__N_2673[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[77] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1429.GSR = "ENABLED";
    FD1P3AX array_255___i1430 (.D(array_0__7__N_2673[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[77] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1430.GSR = "ENABLED";
    FD1P3AX array_255___i1431 (.D(array_0__7__N_2673[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[77] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1431.GSR = "ENABLED";
    FD1P3AX array_255___i1432 (.D(array_0__7__N_2673[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[77] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1432.GSR = "ENABLED";
    FD1P3AX array_255___i1433 (.D(array_0__7__N_2665[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[76] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1433.GSR = "ENABLED";
    FD1P3AX array_255___i1434 (.D(array_0__7__N_2665[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[76] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1434.GSR = "ENABLED";
    FD1P3AX array_255___i1435 (.D(array_0__7__N_2665[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[76] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1435.GSR = "ENABLED";
    FD1P3AX array_255___i1436 (.D(array_0__7__N_2665[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[76] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1436.GSR = "ENABLED";
    FD1P3AX array_255___i1437 (.D(array_0__7__N_2665[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[76] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1437.GSR = "ENABLED";
    FD1P3AX array_255___i1438 (.D(array_0__7__N_2665[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[76] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1438.GSR = "ENABLED";
    FD1P3AX array_255___i1439 (.D(array_0__7__N_2665[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[76] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1439.GSR = "ENABLED";
    FD1P3AX array_255___i1440 (.D(array_0__7__N_2665[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[76] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1440.GSR = "ENABLED";
    FD1P3AX array_255___i1441 (.D(array_0__7__N_2657[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[75] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1441.GSR = "ENABLED";
    FD1P3AX array_255___i1442 (.D(array_0__7__N_2657[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[75] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1442.GSR = "ENABLED";
    FD1P3AX array_255___i1443 (.D(array_0__7__N_2657[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[75] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1443.GSR = "ENABLED";
    FD1P3AX array_255___i1444 (.D(array_0__7__N_2657[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[75] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1444.GSR = "ENABLED";
    FD1P3AX array_255___i1445 (.D(array_0__7__N_2657[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[75] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1445.GSR = "ENABLED";
    FD1P3AX array_255___i1446 (.D(array_0__7__N_2657[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[75] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1446.GSR = "ENABLED";
    FD1P3AX array_255___i1447 (.D(array_0__7__N_2657[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[75] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1447.GSR = "ENABLED";
    FD1P3AX array_255___i1448 (.D(array_0__7__N_2657[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[75] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1448.GSR = "ENABLED";
    FD1P3AX array_255___i1449 (.D(array_0__7__N_2649[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[74] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1449.GSR = "ENABLED";
    FD1P3AX array_255___i1450 (.D(array_0__7__N_2649[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[74] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1450.GSR = "ENABLED";
    FD1P3AX array_255___i1451 (.D(array_0__7__N_2649[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[74] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1451.GSR = "ENABLED";
    FD1P3AX array_255___i1452 (.D(array_0__7__N_2649[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[74] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1452.GSR = "ENABLED";
    FD1P3AX array_255___i1453 (.D(array_0__7__N_2649[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[74] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1453.GSR = "ENABLED";
    FD1P3AX array_255___i1454 (.D(array_0__7__N_2649[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[74] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1454.GSR = "ENABLED";
    FD1P3AX array_255___i1455 (.D(array_0__7__N_2649[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[74] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1455.GSR = "ENABLED";
    FD1P3AX array_255___i1456 (.D(array_0__7__N_2649[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[74] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1456.GSR = "ENABLED";
    FD1P3AX array_255___i1457 (.D(array_0__7__N_2641[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[73] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1457.GSR = "ENABLED";
    FD1P3AX array_255___i1458 (.D(array_0__7__N_2641[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[73] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1458.GSR = "ENABLED";
    FD1P3AX array_255___i1459 (.D(array_0__7__N_2641[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[73] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1459.GSR = "ENABLED";
    FD1P3AX array_255___i1460 (.D(array_0__7__N_2641[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[73] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1460.GSR = "ENABLED";
    FD1P3AX array_255___i1461 (.D(array_0__7__N_2641[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[73] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1461.GSR = "ENABLED";
    FD1P3AX array_255___i1462 (.D(array_0__7__N_2641[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[73] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1462.GSR = "ENABLED";
    FD1P3AX array_255___i1463 (.D(array_0__7__N_2641[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[73] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1463.GSR = "ENABLED";
    FD1P3AX array_255___i1464 (.D(array_0__7__N_2641[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[73] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1464.GSR = "ENABLED";
    FD1P3AX array_255___i1465 (.D(array_0__7__N_2633[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[72] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1465.GSR = "ENABLED";
    FD1P3AX array_255___i1466 (.D(array_0__7__N_2633[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[72] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1466.GSR = "ENABLED";
    FD1P3AX array_255___i1467 (.D(array_0__7__N_2633[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[72] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1467.GSR = "ENABLED";
    FD1P3AX array_255___i1468 (.D(array_0__7__N_2633[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[72] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1468.GSR = "ENABLED";
    FD1P3AX array_255___i1469 (.D(array_0__7__N_2633[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[72] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1469.GSR = "ENABLED";
    FD1P3AX array_255___i1470 (.D(array_0__7__N_2633[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[72] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1470.GSR = "ENABLED";
    FD1P3AX array_255___i1471 (.D(array_0__7__N_2633[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[72] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1471.GSR = "ENABLED";
    FD1P3AX array_255___i1472 (.D(array_0__7__N_2633[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[72] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1472.GSR = "ENABLED";
    FD1P3AX array_255___i1473 (.D(array_0__7__N_2625[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[71] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1473.GSR = "ENABLED";
    FD1P3AX array_255___i1474 (.D(array_0__7__N_2625[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[71] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1474.GSR = "ENABLED";
    FD1P3AX array_255___i1475 (.D(array_0__7__N_2625[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[71] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1475.GSR = "ENABLED";
    FD1P3AX array_255___i1476 (.D(array_0__7__N_2625[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[71] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1476.GSR = "ENABLED";
    FD1P3AX array_255___i1477 (.D(array_0__7__N_2625[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[71] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1477.GSR = "ENABLED";
    FD1P3AX array_255___i1478 (.D(array_0__7__N_2625[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[71] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1478.GSR = "ENABLED";
    FD1P3AX array_255___i1479 (.D(array_0__7__N_2625[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[71] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1479.GSR = "ENABLED";
    FD1P3AX array_255___i1480 (.D(array_0__7__N_2625[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[71] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1480.GSR = "ENABLED";
    FD1P3AX array_255___i1481 (.D(array_0__7__N_2617[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[70] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1481.GSR = "ENABLED";
    FD1P3AX array_255___i1482 (.D(array_0__7__N_2617[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[70] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1482.GSR = "ENABLED";
    FD1P3AX array_255___i1483 (.D(array_0__7__N_2617[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[70] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1483.GSR = "ENABLED";
    FD1P3AX array_255___i1484 (.D(array_0__7__N_2617[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[70] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1484.GSR = "ENABLED";
    FD1P3AX array_255___i1485 (.D(array_0__7__N_2617[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[70] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1485.GSR = "ENABLED";
    FD1P3AX array_255___i1486 (.D(array_0__7__N_2617[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[70] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1486.GSR = "ENABLED";
    FD1P3AX array_255___i1487 (.D(array_0__7__N_2617[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[70] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1487.GSR = "ENABLED";
    FD1P3AX array_255___i1488 (.D(array_0__7__N_2617[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[70] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1488.GSR = "ENABLED";
    FD1P3AX array_255___i1489 (.D(array_0__7__N_2609[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[69] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1489.GSR = "ENABLED";
    FD1P3AX array_255___i1490 (.D(array_0__7__N_2609[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[69] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1490.GSR = "ENABLED";
    FD1P3AX array_255___i1491 (.D(array_0__7__N_2609[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[69] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1491.GSR = "ENABLED";
    FD1P3AX array_255___i1492 (.D(array_0__7__N_2609[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[69] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1492.GSR = "ENABLED";
    FD1P3AX array_255___i1493 (.D(array_0__7__N_2609[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[69] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1493.GSR = "ENABLED";
    FD1P3AX array_255___i1494 (.D(array_0__7__N_2609[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[69] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1494.GSR = "ENABLED";
    FD1P3AX array_255___i1495 (.D(array_0__7__N_2609[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[69] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1495.GSR = "ENABLED";
    FD1P3AX array_255___i1496 (.D(array_0__7__N_2609[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[69] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1496.GSR = "ENABLED";
    FD1P3AX array_255___i1497 (.D(array_0__7__N_2601[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[68] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1497.GSR = "ENABLED";
    FD1P3AX array_255___i1498 (.D(array_0__7__N_2601[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[68] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1498.GSR = "ENABLED";
    FD1P3AX array_255___i1499 (.D(array_0__7__N_2601[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[68] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1499.GSR = "ENABLED";
    FD1P3AX array_255___i1500 (.D(array_0__7__N_2601[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[68] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1500.GSR = "ENABLED";
    FD1P3AX array_255___i1501 (.D(array_0__7__N_2601[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[68] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1501.GSR = "ENABLED";
    FD1P3AX array_255___i1502 (.D(array_0__7__N_2601[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[68] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1502.GSR = "ENABLED";
    FD1P3AX array_255___i1503 (.D(array_0__7__N_2601[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[68] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1503.GSR = "ENABLED";
    FD1P3AX array_255___i1504 (.D(array_0__7__N_2601[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[68] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1504.GSR = "ENABLED";
    FD1P3AX array_255___i1505 (.D(array_0__7__N_2593[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[67] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1505.GSR = "ENABLED";
    FD1P3AX array_255___i1506 (.D(array_0__7__N_2593[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[67] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1506.GSR = "ENABLED";
    FD1P3AX array_255___i1507 (.D(array_0__7__N_2593[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[67] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1507.GSR = "ENABLED";
    FD1P3AX array_255___i1508 (.D(array_0__7__N_2593[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[67] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1508.GSR = "ENABLED";
    FD1P3AX array_255___i1509 (.D(array_0__7__N_2593[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[67] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1509.GSR = "ENABLED";
    FD1P3AX array_255___i1510 (.D(array_0__7__N_2593[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[67] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1510.GSR = "ENABLED";
    FD1P3AX array_255___i1511 (.D(array_0__7__N_2593[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[67] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1511.GSR = "ENABLED";
    FD1P3AX array_255___i1512 (.D(array_0__7__N_2593[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[67] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1512.GSR = "ENABLED";
    FD1P3AX array_255___i1513 (.D(array_0__7__N_2585[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[66] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1513.GSR = "ENABLED";
    FD1P3AX array_255___i1514 (.D(array_0__7__N_2585[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[66] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1514.GSR = "ENABLED";
    FD1P3AX array_255___i1515 (.D(array_0__7__N_2585[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[66] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1515.GSR = "ENABLED";
    FD1P3AX array_255___i1516 (.D(array_0__7__N_2585[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[66] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1516.GSR = "ENABLED";
    FD1P3AX array_255___i1517 (.D(array_0__7__N_2585[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[66] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1517.GSR = "ENABLED";
    FD1P3AX array_255___i1518 (.D(array_0__7__N_2585[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[66] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1518.GSR = "ENABLED";
    FD1P3AX array_255___i1519 (.D(array_0__7__N_2585[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[66] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1519.GSR = "ENABLED";
    FD1P3AX array_255___i1520 (.D(array_0__7__N_2585[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[66] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1520.GSR = "ENABLED";
    FD1P3AX array_255___i1521 (.D(array_0__7__N_2577[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[65] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1521.GSR = "ENABLED";
    FD1P3AX array_255___i1522 (.D(array_0__7__N_2577[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[65] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1522.GSR = "ENABLED";
    FD1P3AX array_255___i1523 (.D(array_0__7__N_2577[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[65] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1523.GSR = "ENABLED";
    FD1P3AX array_255___i1524 (.D(array_0__7__N_2577[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[65] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1524.GSR = "ENABLED";
    FD1P3AX array_255___i1525 (.D(array_0__7__N_2577[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[65] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1525.GSR = "ENABLED";
    FD1P3AX array_255___i1526 (.D(array_0__7__N_2577[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[65] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1526.GSR = "ENABLED";
    FD1P3AX array_255___i1527 (.D(array_0__7__N_2577[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[65] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1527.GSR = "ENABLED";
    FD1P3AX array_255___i1528 (.D(array_0__7__N_2577[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[65] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1528.GSR = "ENABLED";
    FD1P3AX array_255___i1529 (.D(array_0__7__N_2569[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[64] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1529.GSR = "ENABLED";
    FD1P3AX array_255___i1530 (.D(array_0__7__N_2569[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[64] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1530.GSR = "ENABLED";
    FD1P3AX array_255___i1531 (.D(array_0__7__N_2569[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[64] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1531.GSR = "ENABLED";
    FD1P3AX array_255___i1532 (.D(array_0__7__N_2569[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[64] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1532.GSR = "ENABLED";
    FD1P3AX array_255___i1533 (.D(array_0__7__N_2569[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[64] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1533.GSR = "ENABLED";
    FD1P3AX array_255___i1534 (.D(array_0__7__N_2569[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[64] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1534.GSR = "ENABLED";
    FD1P3AX array_255___i1535 (.D(array_0__7__N_2569[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[64] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1535.GSR = "ENABLED";
    FD1P3AX array_255___i1536 (.D(array_0__7__N_2569[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[64] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1536.GSR = "ENABLED";
    FD1P3AX array_255___i1537 (.D(array_0__7__N_2561[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[63] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1537.GSR = "ENABLED";
    FD1P3AX array_255___i1538 (.D(array_0__7__N_2561[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[63] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1538.GSR = "ENABLED";
    FD1P3AX array_255___i1539 (.D(array_0__7__N_2561[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[63] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1539.GSR = "ENABLED";
    FD1P3AX array_255___i1540 (.D(array_0__7__N_2561[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[63] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1540.GSR = "ENABLED";
    FD1P3AX array_255___i1541 (.D(array_0__7__N_2561[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[63] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1541.GSR = "ENABLED";
    FD1P3AX array_255___i1542 (.D(array_0__7__N_2561[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[63] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1542.GSR = "ENABLED";
    FD1P3AX array_255___i1543 (.D(array_0__7__N_2561[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[63] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1543.GSR = "ENABLED";
    FD1P3AX array_255___i1544 (.D(array_0__7__N_2561[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[63] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1544.GSR = "ENABLED";
    FD1P3AX array_255___i1545 (.D(array_0__7__N_2553[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[62] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1545.GSR = "ENABLED";
    FD1P3AX array_255___i1546 (.D(array_0__7__N_2553[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[62] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1546.GSR = "ENABLED";
    FD1P3AX array_255___i1547 (.D(array_0__7__N_2553[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[62] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1547.GSR = "ENABLED";
    FD1P3AX array_255___i1548 (.D(array_0__7__N_2553[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[62] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1548.GSR = "ENABLED";
    FD1P3AX array_255___i1549 (.D(array_0__7__N_2553[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[62] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1549.GSR = "ENABLED";
    FD1P3AX array_255___i1550 (.D(array_0__7__N_2553[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[62] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1550.GSR = "ENABLED";
    FD1P3AX array_255___i1551 (.D(array_0__7__N_2553[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[62] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1551.GSR = "ENABLED";
    FD1P3AX array_255___i1552 (.D(array_0__7__N_2553[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[62] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1552.GSR = "ENABLED";
    FD1P3AX array_255___i1553 (.D(array_0__7__N_2545[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[61] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1553.GSR = "ENABLED";
    FD1P3AX array_255___i1554 (.D(array_0__7__N_2545[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[61] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1554.GSR = "ENABLED";
    FD1P3AX array_255___i1555 (.D(array_0__7__N_2545[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[61] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1555.GSR = "ENABLED";
    FD1P3AX array_255___i1556 (.D(array_0__7__N_2545[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[61] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1556.GSR = "ENABLED";
    FD1P3AX array_255___i1557 (.D(array_0__7__N_2545[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[61] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1557.GSR = "ENABLED";
    FD1P3AX array_255___i1558 (.D(array_0__7__N_2545[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[61] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1558.GSR = "ENABLED";
    FD1P3AX array_255___i1559 (.D(array_0__7__N_2545[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[61] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1559.GSR = "ENABLED";
    FD1P3AX array_255___i1560 (.D(array_0__7__N_2545[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[61] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1560.GSR = "ENABLED";
    FD1P3AX array_255___i1561 (.D(array_0__7__N_2537[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[60] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1561.GSR = "ENABLED";
    FD1P3AX array_255___i1562 (.D(array_0__7__N_2537[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[60] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1562.GSR = "ENABLED";
    FD1P3AX array_255___i1563 (.D(array_0__7__N_2537[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[60] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1563.GSR = "ENABLED";
    FD1P3AX array_255___i1564 (.D(array_0__7__N_2537[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[60] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1564.GSR = "ENABLED";
    FD1P3AX array_255___i1565 (.D(array_0__7__N_2537[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[60] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1565.GSR = "ENABLED";
    FD1P3AX array_255___i1566 (.D(array_0__7__N_2537[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[60] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1566.GSR = "ENABLED";
    FD1P3AX array_255___i1567 (.D(array_0__7__N_2537[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[60] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1567.GSR = "ENABLED";
    FD1P3AX array_255___i1568 (.D(array_0__7__N_2537[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[60] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1568.GSR = "ENABLED";
    FD1P3AX array_255___i1569 (.D(array_0__7__N_2529[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[59] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1569.GSR = "ENABLED";
    FD1P3AX array_255___i1570 (.D(array_0__7__N_2529[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[59] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1570.GSR = "ENABLED";
    FD1P3AX array_255___i1571 (.D(array_0__7__N_2529[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[59] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1571.GSR = "ENABLED";
    FD1P3AX array_255___i1572 (.D(array_0__7__N_2529[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[59] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1572.GSR = "ENABLED";
    FD1P3AX array_255___i1573 (.D(array_0__7__N_2529[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[59] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1573.GSR = "ENABLED";
    FD1P3AX array_255___i1574 (.D(array_0__7__N_2529[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[59] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1574.GSR = "ENABLED";
    FD1P3AX array_255___i1575 (.D(array_0__7__N_2529[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[59] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1575.GSR = "ENABLED";
    FD1P3AX array_255___i1576 (.D(array_0__7__N_2529[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[59] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1576.GSR = "ENABLED";
    FD1P3AX array_255___i1577 (.D(array_0__7__N_2521[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[58] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1577.GSR = "ENABLED";
    FD1P3AX array_255___i1578 (.D(array_0__7__N_2521[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[58] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1578.GSR = "ENABLED";
    FD1P3AX array_255___i1579 (.D(array_0__7__N_2521[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[58] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1579.GSR = "ENABLED";
    FD1P3AX array_255___i1580 (.D(array_0__7__N_2521[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[58] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1580.GSR = "ENABLED";
    FD1P3AX array_255___i1581 (.D(array_0__7__N_2521[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[58] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1581.GSR = "ENABLED";
    FD1P3AX array_255___i1582 (.D(array_0__7__N_2521[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[58] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1582.GSR = "ENABLED";
    FD1P3AX array_255___i1583 (.D(array_0__7__N_2521[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[58] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1583.GSR = "ENABLED";
    FD1P3AX array_255___i1584 (.D(array_0__7__N_2521[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[58] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1584.GSR = "ENABLED";
    FD1P3AX array_255___i1585 (.D(array_0__7__N_2513[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[57] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1585.GSR = "ENABLED";
    FD1P3AX array_255___i1586 (.D(array_0__7__N_2513[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[57] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1586.GSR = "ENABLED";
    FD1P3AX array_255___i1587 (.D(array_0__7__N_2513[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[57] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1587.GSR = "ENABLED";
    FD1P3AX array_255___i1588 (.D(array_0__7__N_2513[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[57] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1588.GSR = "ENABLED";
    FD1P3AX array_255___i1589 (.D(array_0__7__N_2513[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[57] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1589.GSR = "ENABLED";
    FD1P3AX array_255___i1590 (.D(array_0__7__N_2513[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[57] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1590.GSR = "ENABLED";
    FD1P3AX array_255___i1591 (.D(array_0__7__N_2513[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[57] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1591.GSR = "ENABLED";
    FD1P3AX array_255___i1592 (.D(array_0__7__N_2513[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[57] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1592.GSR = "ENABLED";
    FD1P3AX array_255___i1593 (.D(array_0__7__N_2505[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[56] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1593.GSR = "ENABLED";
    FD1P3AX array_255___i1594 (.D(array_0__7__N_2505[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[56] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1594.GSR = "ENABLED";
    FD1P3AX array_255___i1595 (.D(array_0__7__N_2505[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[56] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1595.GSR = "ENABLED";
    FD1P3AX array_255___i1596 (.D(array_0__7__N_2505[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[56] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1596.GSR = "ENABLED";
    FD1P3AX array_255___i1597 (.D(array_0__7__N_2505[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[56] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1597.GSR = "ENABLED";
    FD1P3AX array_255___i1598 (.D(array_0__7__N_2505[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[56] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1598.GSR = "ENABLED";
    FD1P3AX array_255___i1599 (.D(array_0__7__N_2505[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[56] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1599.GSR = "ENABLED";
    FD1P3AX array_255___i1600 (.D(array_0__7__N_2505[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[56] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1600.GSR = "ENABLED";
    FD1P3AX array_255___i1601 (.D(array_0__7__N_2497[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[55] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1601.GSR = "ENABLED";
    FD1P3AX array_255___i1602 (.D(array_0__7__N_2497[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[55] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1602.GSR = "ENABLED";
    FD1P3AX array_255___i1603 (.D(array_0__7__N_2497[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[55] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1603.GSR = "ENABLED";
    FD1P3AX array_255___i1604 (.D(array_0__7__N_2497[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[55] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1604.GSR = "ENABLED";
    FD1P3AX array_255___i1605 (.D(array_0__7__N_2497[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[55] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1605.GSR = "ENABLED";
    FD1P3AX array_255___i1606 (.D(array_0__7__N_2497[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[55] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1606.GSR = "ENABLED";
    FD1P3AX array_255___i1607 (.D(array_0__7__N_2497[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[55] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1607.GSR = "ENABLED";
    FD1P3AX array_255___i1608 (.D(array_0__7__N_2497[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[55] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1608.GSR = "ENABLED";
    FD1P3AX array_255___i1609 (.D(array_0__7__N_2489[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[54] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1609.GSR = "ENABLED";
    FD1P3AX array_255___i1610 (.D(array_0__7__N_2489[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[54] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1610.GSR = "ENABLED";
    FD1P3AX array_255___i1611 (.D(array_0__7__N_2489[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[54] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1611.GSR = "ENABLED";
    FD1P3AX array_255___i1612 (.D(array_0__7__N_2489[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[54] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1612.GSR = "ENABLED";
    FD1P3AX array_255___i1613 (.D(array_0__7__N_2489[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[54] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1613.GSR = "ENABLED";
    FD1P3AX array_255___i1614 (.D(array_0__7__N_2489[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[54] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1614.GSR = "ENABLED";
    FD1P3AX array_255___i1615 (.D(array_0__7__N_2489[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[54] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1615.GSR = "ENABLED";
    FD1P3AX array_255___i1616 (.D(array_0__7__N_2489[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[54] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1616.GSR = "ENABLED";
    FD1P3AX array_255___i1617 (.D(array_0__7__N_2481[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[53] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1617.GSR = "ENABLED";
    FD1P3AX array_255___i1618 (.D(array_0__7__N_2481[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[53] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1618.GSR = "ENABLED";
    FD1P3AX array_255___i1619 (.D(array_0__7__N_2481[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[53] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1619.GSR = "ENABLED";
    FD1P3AX array_255___i1620 (.D(array_0__7__N_2481[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[53] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1620.GSR = "ENABLED";
    FD1P3AX array_255___i1621 (.D(array_0__7__N_2481[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[53] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1621.GSR = "ENABLED";
    FD1P3AX array_255___i1622 (.D(array_0__7__N_2481[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[53] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1622.GSR = "ENABLED";
    FD1P3AX array_255___i1623 (.D(array_0__7__N_2481[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[53] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1623.GSR = "ENABLED";
    FD1P3AX array_255___i1624 (.D(array_0__7__N_2481[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[53] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1624.GSR = "ENABLED";
    FD1P3AX array_255___i1625 (.D(array_0__7__N_2473[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[52] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1625.GSR = "ENABLED";
    FD1P3AX array_255___i1626 (.D(array_0__7__N_2473[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[52] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1626.GSR = "ENABLED";
    FD1P3AX array_255___i1627 (.D(array_0__7__N_2473[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[52] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1627.GSR = "ENABLED";
    FD1P3AX array_255___i1628 (.D(array_0__7__N_2473[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[52] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1628.GSR = "ENABLED";
    FD1P3AX array_255___i1629 (.D(array_0__7__N_2473[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[52] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1629.GSR = "ENABLED";
    FD1P3AX array_255___i1630 (.D(array_0__7__N_2473[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[52] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1630.GSR = "ENABLED";
    FD1P3AX array_255___i1631 (.D(array_0__7__N_2473[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[52] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1631.GSR = "ENABLED";
    FD1P3AX array_255___i1632 (.D(array_0__7__N_2473[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[52] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1632.GSR = "ENABLED";
    FD1P3AX array_255___i1633 (.D(array_0__7__N_2465[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[51] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1633.GSR = "ENABLED";
    FD1P3AX array_255___i1634 (.D(array_0__7__N_2465[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[51] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1634.GSR = "ENABLED";
    FD1P3AX array_255___i1635 (.D(array_0__7__N_2465[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[51] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1635.GSR = "ENABLED";
    FD1P3AX array_255___i1636 (.D(array_0__7__N_2465[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[51] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1636.GSR = "ENABLED";
    FD1P3AX array_255___i1637 (.D(array_0__7__N_2465[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[51] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1637.GSR = "ENABLED";
    FD1P3AX array_255___i1638 (.D(array_0__7__N_2465[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[51] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1638.GSR = "ENABLED";
    FD1P3AX array_255___i1639 (.D(array_0__7__N_2465[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[51] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1639.GSR = "ENABLED";
    FD1P3AX array_255___i1640 (.D(array_0__7__N_2465[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[51] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1640.GSR = "ENABLED";
    FD1P3AX array_255___i1641 (.D(array_0__7__N_2457[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[50] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1641.GSR = "ENABLED";
    FD1P3AX array_255___i1642 (.D(array_0__7__N_2457[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[50] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1642.GSR = "ENABLED";
    FD1P3AX array_255___i1643 (.D(array_0__7__N_2457[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[50] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1643.GSR = "ENABLED";
    FD1P3AX array_255___i1644 (.D(array_0__7__N_2457[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[50] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1644.GSR = "ENABLED";
    FD1P3AX array_255___i1645 (.D(array_0__7__N_2457[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[50] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1645.GSR = "ENABLED";
    FD1P3AX array_255___i1646 (.D(array_0__7__N_2457[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[50] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1646.GSR = "ENABLED";
    FD1P3AX array_255___i1647 (.D(array_0__7__N_2457[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[50] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1647.GSR = "ENABLED";
    FD1P3AX array_255___i1648 (.D(array_0__7__N_2457[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[50] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1648.GSR = "ENABLED";
    FD1P3AX array_255___i1649 (.D(array_0__7__N_2449[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[49] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1649.GSR = "ENABLED";
    FD1P3AX array_255___i1650 (.D(array_0__7__N_2449[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[49] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1650.GSR = "ENABLED";
    FD1P3AX array_255___i1651 (.D(array_0__7__N_2449[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[49] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1651.GSR = "ENABLED";
    FD1P3AX array_255___i1652 (.D(array_0__7__N_2449[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[49] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1652.GSR = "ENABLED";
    FD1P3AX array_255___i1653 (.D(array_0__7__N_2449[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[49] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1653.GSR = "ENABLED";
    FD1P3AX array_255___i1654 (.D(array_0__7__N_2449[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[49] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1654.GSR = "ENABLED";
    FD1P3AX array_255___i1655 (.D(array_0__7__N_2449[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[49] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1655.GSR = "ENABLED";
    FD1P3AX array_255___i1656 (.D(array_0__7__N_2449[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[49] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1656.GSR = "ENABLED";
    FD1P3AX array_255___i1657 (.D(array_0__7__N_2441[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[48] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1657.GSR = "ENABLED";
    FD1P3AX array_255___i1658 (.D(array_0__7__N_2441[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[48] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1658.GSR = "ENABLED";
    FD1P3AX array_255___i1659 (.D(array_0__7__N_2441[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[48] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1659.GSR = "ENABLED";
    FD1P3AX array_255___i1660 (.D(array_0__7__N_2441[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[48] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1660.GSR = "ENABLED";
    FD1P3AX array_255___i1661 (.D(array_0__7__N_2441[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[48] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1661.GSR = "ENABLED";
    FD1P3AX array_255___i1662 (.D(array_0__7__N_2441[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[48] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1662.GSR = "ENABLED";
    FD1P3AX array_255___i1663 (.D(array_0__7__N_2441[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[48] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1663.GSR = "ENABLED";
    FD1P3AX array_255___i1664 (.D(array_0__7__N_2441[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[48] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1664.GSR = "ENABLED";
    FD1P3AX array_255___i1665 (.D(array_0__7__N_2433[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[47] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1665.GSR = "ENABLED";
    FD1P3AX array_255___i1666 (.D(array_0__7__N_2433[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[47] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1666.GSR = "ENABLED";
    FD1P3AX array_255___i1667 (.D(array_0__7__N_2433[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[47] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1667.GSR = "ENABLED";
    FD1P3AX array_255___i1668 (.D(array_0__7__N_2433[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[47] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1668.GSR = "ENABLED";
    FD1P3AX array_255___i1669 (.D(array_0__7__N_2433[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[47] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1669.GSR = "ENABLED";
    FD1P3AX array_255___i1670 (.D(array_0__7__N_2433[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[47] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1670.GSR = "ENABLED";
    FD1P3AX array_255___i1671 (.D(array_0__7__N_2433[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[47] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1671.GSR = "ENABLED";
    FD1P3AX array_255___i1672 (.D(array_0__7__N_2433[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[47] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1672.GSR = "ENABLED";
    FD1P3AX array_255___i1673 (.D(array_0__7__N_2425[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[46] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1673.GSR = "ENABLED";
    FD1P3AX array_255___i1674 (.D(array_0__7__N_2425[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[46] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1674.GSR = "ENABLED";
    FD1P3AX array_255___i1675 (.D(array_0__7__N_2425[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[46] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1675.GSR = "ENABLED";
    FD1P3AX array_255___i1676 (.D(array_0__7__N_2425[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[46] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1676.GSR = "ENABLED";
    FD1P3AX array_255___i1677 (.D(array_0__7__N_2425[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[46] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1677.GSR = "ENABLED";
    FD1P3AX array_255___i1678 (.D(array_0__7__N_2425[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[46] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1678.GSR = "ENABLED";
    FD1P3AX array_255___i1679 (.D(array_0__7__N_2425[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[46] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1679.GSR = "ENABLED";
    FD1P3AX array_255___i1680 (.D(array_0__7__N_2425[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[46] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1680.GSR = "ENABLED";
    FD1P3AX array_255___i1681 (.D(array_0__7__N_2417[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[45] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1681.GSR = "ENABLED";
    FD1P3AX array_255___i1682 (.D(array_0__7__N_2417[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[45] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1682.GSR = "ENABLED";
    FD1P3AX array_255___i1683 (.D(array_0__7__N_2417[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[45] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1683.GSR = "ENABLED";
    FD1P3AX array_255___i1684 (.D(array_0__7__N_2417[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[45] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1684.GSR = "ENABLED";
    FD1P3AX array_255___i1685 (.D(array_0__7__N_2417[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[45] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1685.GSR = "ENABLED";
    FD1P3AX array_255___i1686 (.D(array_0__7__N_2417[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[45] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1686.GSR = "ENABLED";
    FD1P3AX array_255___i1687 (.D(array_0__7__N_2417[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[45] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1687.GSR = "ENABLED";
    FD1P3AX array_255___i1688 (.D(array_0__7__N_2417[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[45] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1688.GSR = "ENABLED";
    FD1P3AX array_255___i1689 (.D(array_0__7__N_2409[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[44] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1689.GSR = "ENABLED";
    FD1P3AX array_255___i1690 (.D(array_0__7__N_2409[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[44] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1690.GSR = "ENABLED";
    FD1P3AX array_255___i1691 (.D(array_0__7__N_2409[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[44] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1691.GSR = "ENABLED";
    FD1P3AX array_255___i1692 (.D(array_0__7__N_2409[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[44] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1692.GSR = "ENABLED";
    FD1P3AX array_255___i1693 (.D(array_0__7__N_2409[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[44] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1693.GSR = "ENABLED";
    FD1P3AX array_255___i1694 (.D(array_0__7__N_2409[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[44] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1694.GSR = "ENABLED";
    FD1P3AX array_255___i1695 (.D(array_0__7__N_2409[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[44] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1695.GSR = "ENABLED";
    FD1P3AX array_255___i1696 (.D(array_0__7__N_2409[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[44] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1696.GSR = "ENABLED";
    FD1P3AX array_255___i1697 (.D(array_0__7__N_2401[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[43] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1697.GSR = "ENABLED";
    FD1P3AX array_255___i1698 (.D(array_0__7__N_2401[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[43] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1698.GSR = "ENABLED";
    FD1P3AX array_255___i1699 (.D(array_0__7__N_2401[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[43] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1699.GSR = "ENABLED";
    FD1P3AX array_255___i1700 (.D(array_0__7__N_2401[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[43] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1700.GSR = "ENABLED";
    FD1P3AX array_255___i1701 (.D(array_0__7__N_2401[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[43] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1701.GSR = "ENABLED";
    FD1P3AX array_255___i1702 (.D(array_0__7__N_2401[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[43] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1702.GSR = "ENABLED";
    FD1P3AX array_255___i1703 (.D(array_0__7__N_2401[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[43] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1703.GSR = "ENABLED";
    FD1P3AX array_255___i1704 (.D(array_0__7__N_2401[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[43] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1704.GSR = "ENABLED";
    FD1P3AX array_255___i1705 (.D(array_0__7__N_2393[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[42] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1705.GSR = "ENABLED";
    FD1P3AX array_255___i1706 (.D(array_0__7__N_2393[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[42] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1706.GSR = "ENABLED";
    FD1P3AX array_255___i1707 (.D(array_0__7__N_2393[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[42] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1707.GSR = "ENABLED";
    FD1P3AX array_255___i1708 (.D(array_0__7__N_2393[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[42] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1708.GSR = "ENABLED";
    FD1P3AX array_255___i1709 (.D(array_0__7__N_2393[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[42] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1709.GSR = "ENABLED";
    FD1P3AX array_255___i1710 (.D(array_0__7__N_2393[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[42] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1710.GSR = "ENABLED";
    FD1P3AX array_255___i1711 (.D(array_0__7__N_2393[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[42] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1711.GSR = "ENABLED";
    FD1P3AX array_255___i1712 (.D(array_0__7__N_2393[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[42] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1712.GSR = "ENABLED";
    FD1P3AX array_255___i1713 (.D(array_0__7__N_2385[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[41] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1713.GSR = "ENABLED";
    FD1P3AX array_255___i1714 (.D(array_0__7__N_2385[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[41] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1714.GSR = "ENABLED";
    FD1P3AX array_255___i1715 (.D(array_0__7__N_2385[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[41] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1715.GSR = "ENABLED";
    FD1P3AX array_255___i1716 (.D(array_0__7__N_2385[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[41] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1716.GSR = "ENABLED";
    FD1P3AX array_255___i1717 (.D(array_0__7__N_2385[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[41] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1717.GSR = "ENABLED";
    FD1P3AX array_255___i1718 (.D(array_0__7__N_2385[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[41] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1718.GSR = "ENABLED";
    FD1P3AX array_255___i1719 (.D(array_0__7__N_2385[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[41] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1719.GSR = "ENABLED";
    FD1P3AX array_255___i1720 (.D(array_0__7__N_2385[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[41] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1720.GSR = "ENABLED";
    FD1P3AX array_255___i1721 (.D(array_0__7__N_2377[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[40] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1721.GSR = "ENABLED";
    FD1P3AX array_255___i1722 (.D(array_0__7__N_2377[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[40] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1722.GSR = "ENABLED";
    FD1P3AX array_255___i1723 (.D(array_0__7__N_2377[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[40] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1723.GSR = "ENABLED";
    FD1P3AX array_255___i1724 (.D(array_0__7__N_2377[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[40] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1724.GSR = "ENABLED";
    FD1P3AX array_255___i1725 (.D(array_0__7__N_2377[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[40] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1725.GSR = "ENABLED";
    FD1P3AX array_255___i1726 (.D(array_0__7__N_2377[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[40] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1726.GSR = "ENABLED";
    FD1P3AX array_255___i1727 (.D(array_0__7__N_2377[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[40] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1727.GSR = "ENABLED";
    FD1P3AX array_255___i1728 (.D(array_0__7__N_2377[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[40] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1728.GSR = "ENABLED";
    FD1P3AX array_255___i1729 (.D(array_0__7__N_2369[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[39] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1729.GSR = "ENABLED";
    FD1P3AX array_255___i1730 (.D(array_0__7__N_2369[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[39] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1730.GSR = "ENABLED";
    FD1P3AX array_255___i1731 (.D(array_0__7__N_2369[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[39] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1731.GSR = "ENABLED";
    FD1P3AX array_255___i1732 (.D(array_0__7__N_2369[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[39] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1732.GSR = "ENABLED";
    FD1P3AX array_255___i1733 (.D(array_0__7__N_2369[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[39] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1733.GSR = "ENABLED";
    FD1P3AX array_255___i1734 (.D(array_0__7__N_2369[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[39] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1734.GSR = "ENABLED";
    FD1P3AX array_255___i1735 (.D(array_0__7__N_2369[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[39] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1735.GSR = "ENABLED";
    FD1P3AX array_255___i1736 (.D(array_0__7__N_2369[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[39] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1736.GSR = "ENABLED";
    FD1P3AX array_255___i1737 (.D(array_0__7__N_2361[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[38] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1737.GSR = "ENABLED";
    FD1P3AX array_255___i1738 (.D(array_0__7__N_2361[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[38] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1738.GSR = "ENABLED";
    FD1P3AX array_255___i1739 (.D(array_0__7__N_2361[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[38] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1739.GSR = "ENABLED";
    FD1P3AX array_255___i1740 (.D(array_0__7__N_2361[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[38] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1740.GSR = "ENABLED";
    FD1P3AX array_255___i1741 (.D(array_0__7__N_2361[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[38] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1741.GSR = "ENABLED";
    FD1P3AX array_255___i1742 (.D(array_0__7__N_2361[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[38] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1742.GSR = "ENABLED";
    FD1P3AX array_255___i1743 (.D(array_0__7__N_2361[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[38] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1743.GSR = "ENABLED";
    FD1P3AX array_255___i1744 (.D(array_0__7__N_2361[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[38] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1744.GSR = "ENABLED";
    FD1P3AX array_255___i1745 (.D(array_0__7__N_2353[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[37] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1745.GSR = "ENABLED";
    FD1P3AX array_255___i1746 (.D(array_0__7__N_2353[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[37] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1746.GSR = "ENABLED";
    FD1P3AX array_255___i1747 (.D(array_0__7__N_2353[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[37] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1747.GSR = "ENABLED";
    FD1P3AX array_255___i1748 (.D(array_0__7__N_2353[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[37] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1748.GSR = "ENABLED";
    FD1P3AX array_255___i1749 (.D(array_0__7__N_2353[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[37] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1749.GSR = "ENABLED";
    FD1P3AX array_255___i1750 (.D(array_0__7__N_2353[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[37] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1750.GSR = "ENABLED";
    FD1P3AX array_255___i1751 (.D(array_0__7__N_2353[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[37] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1751.GSR = "ENABLED";
    FD1P3AX array_255___i1752 (.D(array_0__7__N_2353[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[37] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1752.GSR = "ENABLED";
    FD1P3AX array_255___i1753 (.D(array_0__7__N_2345[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[36] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1753.GSR = "ENABLED";
    FD1P3AX array_255___i1754 (.D(array_0__7__N_2345[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[36] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1754.GSR = "ENABLED";
    FD1P3AX array_255___i1755 (.D(array_0__7__N_2345[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[36] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1755.GSR = "ENABLED";
    FD1P3AX array_255___i1756 (.D(array_0__7__N_2345[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[36] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1756.GSR = "ENABLED";
    FD1P3AX array_255___i1757 (.D(array_0__7__N_2345[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[36] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1757.GSR = "ENABLED";
    FD1P3AX array_255___i1758 (.D(array_0__7__N_2345[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[36] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1758.GSR = "ENABLED";
    FD1P3AX array_255___i1759 (.D(array_0__7__N_2345[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[36] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1759.GSR = "ENABLED";
    FD1P3AX array_255___i1760 (.D(array_0__7__N_2345[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[36] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1760.GSR = "ENABLED";
    FD1P3AX array_255___i1761 (.D(array_0__7__N_2337[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[35] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1761.GSR = "ENABLED";
    FD1P3AX array_255___i1762 (.D(array_0__7__N_2337[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[35] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1762.GSR = "ENABLED";
    FD1P3AX array_255___i1763 (.D(array_0__7__N_2337[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[35] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1763.GSR = "ENABLED";
    FD1P3AX array_255___i1764 (.D(array_0__7__N_2337[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[35] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1764.GSR = "ENABLED";
    FD1P3AX array_255___i1765 (.D(array_0__7__N_2337[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[35] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1765.GSR = "ENABLED";
    FD1P3AX array_255___i1766 (.D(array_0__7__N_2337[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[35] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1766.GSR = "ENABLED";
    FD1P3AX array_255___i1767 (.D(array_0__7__N_2337[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[35] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1767.GSR = "ENABLED";
    FD1P3AX array_255___i1768 (.D(array_0__7__N_2337[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[35] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1768.GSR = "ENABLED";
    FD1P3AX array_255___i1769 (.D(array_0__7__N_2329[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[34] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1769.GSR = "ENABLED";
    FD1P3AX array_255___i1770 (.D(array_0__7__N_2329[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[34] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1770.GSR = "ENABLED";
    FD1P3AX array_255___i1771 (.D(array_0__7__N_2329[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[34] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1771.GSR = "ENABLED";
    FD1P3AX array_255___i1772 (.D(array_0__7__N_2329[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[34] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1772.GSR = "ENABLED";
    FD1P3AX array_255___i1773 (.D(array_0__7__N_2329[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[34] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1773.GSR = "ENABLED";
    FD1P3AX array_255___i1774 (.D(array_0__7__N_2329[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[34] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1774.GSR = "ENABLED";
    FD1P3AX array_255___i1775 (.D(array_0__7__N_2329[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[34] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1775.GSR = "ENABLED";
    FD1P3AX array_255___i1776 (.D(array_0__7__N_2329[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[34] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1776.GSR = "ENABLED";
    FD1P3AX array_255___i1777 (.D(array_0__7__N_2321[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[33] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1777.GSR = "ENABLED";
    FD1P3AX array_255___i1778 (.D(array_0__7__N_2321[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[33] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1778.GSR = "ENABLED";
    FD1P3AX array_255___i1779 (.D(array_0__7__N_2321[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[33] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1779.GSR = "ENABLED";
    FD1P3AX array_255___i1780 (.D(array_0__7__N_2321[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[33] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1780.GSR = "ENABLED";
    FD1P3AX array_255___i1781 (.D(array_0__7__N_2321[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[33] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1781.GSR = "ENABLED";
    FD1P3AX array_255___i1782 (.D(array_0__7__N_2321[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[33] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1782.GSR = "ENABLED";
    FD1P3AX array_255___i1783 (.D(array_0__7__N_2321[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[33] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1783.GSR = "ENABLED";
    FD1P3AX array_255___i1784 (.D(array_0__7__N_2321[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[33] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1784.GSR = "ENABLED";
    FD1P3AX array_255___i1785 (.D(array_0__7__N_2313[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[32] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1785.GSR = "ENABLED";
    FD1P3AX array_255___i1786 (.D(array_0__7__N_2313[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[32] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1786.GSR = "ENABLED";
    FD1P3AX array_255___i1787 (.D(array_0__7__N_2313[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[32] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1787.GSR = "ENABLED";
    FD1P3AX array_255___i1788 (.D(array_0__7__N_2313[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[32] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1788.GSR = "ENABLED";
    FD1P3AX array_255___i1789 (.D(array_0__7__N_2313[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[32] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1789.GSR = "ENABLED";
    FD1P3AX array_255___i1790 (.D(array_0__7__N_2313[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[32] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1790.GSR = "ENABLED";
    FD1P3AX array_255___i1791 (.D(array_0__7__N_2313[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[32] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1791.GSR = "ENABLED";
    FD1P3AX array_255___i1792 (.D(array_0__7__N_2313[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[32] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1792.GSR = "ENABLED";
    FD1P3AX array_255___i1793 (.D(array_0__7__N_2305[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[31] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1793.GSR = "ENABLED";
    FD1P3AX array_255___i1794 (.D(array_0__7__N_2305[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[31] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1794.GSR = "ENABLED";
    FD1P3AX array_255___i1795 (.D(array_0__7__N_2305[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[31] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1795.GSR = "ENABLED";
    FD1P3AX array_255___i1796 (.D(array_0__7__N_2305[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[31] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1796.GSR = "ENABLED";
    FD1P3AX array_255___i1797 (.D(array_0__7__N_2305[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[31] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1797.GSR = "ENABLED";
    FD1P3AX array_255___i1798 (.D(array_0__7__N_2305[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[31] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1798.GSR = "ENABLED";
    FD1P3AX array_255___i1799 (.D(array_0__7__N_2305[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[31] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1799.GSR = "ENABLED";
    FD1P3AX array_255___i1800 (.D(array_0__7__N_2305[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[31] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1800.GSR = "ENABLED";
    FD1P3AX array_255___i1801 (.D(array_0__7__N_2297[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[30] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1801.GSR = "ENABLED";
    FD1P3AX array_255___i1802 (.D(array_0__7__N_2297[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[30] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1802.GSR = "ENABLED";
    FD1P3AX array_255___i1803 (.D(array_0__7__N_2297[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[30] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1803.GSR = "ENABLED";
    FD1P3AX array_255___i1804 (.D(array_0__7__N_2297[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[30] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1804.GSR = "ENABLED";
    FD1P3AX array_255___i1805 (.D(array_0__7__N_2297[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[30] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1805.GSR = "ENABLED";
    FD1P3AX array_255___i1806 (.D(array_0__7__N_2297[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[30] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1806.GSR = "ENABLED";
    FD1P3AX array_255___i1807 (.D(array_0__7__N_2297[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[30] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1807.GSR = "ENABLED";
    FD1P3AX array_255___i1808 (.D(array_0__7__N_2297[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[30] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1808.GSR = "ENABLED";
    FD1P3AX array_255___i1809 (.D(array_0__7__N_2289[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[29] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1809.GSR = "ENABLED";
    FD1P3AX array_255___i1810 (.D(array_0__7__N_2289[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[29] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1810.GSR = "ENABLED";
    FD1P3AX array_255___i1811 (.D(array_0__7__N_2289[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[29] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1811.GSR = "ENABLED";
    FD1P3AX array_255___i1812 (.D(array_0__7__N_2289[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[29] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1812.GSR = "ENABLED";
    FD1P3AX array_255___i1813 (.D(array_0__7__N_2289[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[29] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1813.GSR = "ENABLED";
    FD1P3AX array_255___i1814 (.D(array_0__7__N_2289[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[29] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1814.GSR = "ENABLED";
    FD1P3AX array_255___i1815 (.D(array_0__7__N_2289[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[29] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1815.GSR = "ENABLED";
    FD1P3AX array_255___i1816 (.D(array_0__7__N_2289[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[29] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1816.GSR = "ENABLED";
    FD1P3AX array_255___i1817 (.D(array_0__7__N_2281[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[28] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1817.GSR = "ENABLED";
    FD1P3AX array_255___i1818 (.D(array_0__7__N_2281[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[28] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1818.GSR = "ENABLED";
    FD1P3AX array_255___i1819 (.D(array_0__7__N_2281[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[28] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1819.GSR = "ENABLED";
    FD1P3AX array_255___i1820 (.D(array_0__7__N_2281[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[28] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1820.GSR = "ENABLED";
    FD1P3AX array_255___i1821 (.D(array_0__7__N_2281[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[28] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1821.GSR = "ENABLED";
    FD1P3AX array_255___i1822 (.D(array_0__7__N_2281[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[28] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1822.GSR = "ENABLED";
    FD1P3AX array_255___i1823 (.D(array_0__7__N_2281[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[28] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1823.GSR = "ENABLED";
    FD1P3AX array_255___i1824 (.D(array_0__7__N_2281[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[28] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1824.GSR = "ENABLED";
    FD1P3AX array_255___i1825 (.D(array_0__7__N_2273[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[27] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1825.GSR = "ENABLED";
    FD1P3AX array_255___i1826 (.D(array_0__7__N_2273[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[27] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1826.GSR = "ENABLED";
    FD1P3AX array_255___i1827 (.D(array_0__7__N_2273[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[27] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1827.GSR = "ENABLED";
    FD1P3AX array_255___i1828 (.D(array_0__7__N_2273[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[27] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1828.GSR = "ENABLED";
    FD1P3AX array_255___i1829 (.D(array_0__7__N_2273[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[27] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1829.GSR = "ENABLED";
    FD1P3AX array_255___i1830 (.D(array_0__7__N_2273[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[27] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1830.GSR = "ENABLED";
    FD1P3AX array_255___i1831 (.D(array_0__7__N_2273[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[27] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1831.GSR = "ENABLED";
    FD1P3AX array_255___i1832 (.D(array_0__7__N_2273[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[27] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1832.GSR = "ENABLED";
    FD1P3AX array_255___i1833 (.D(array_0__7__N_2265[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[26] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1833.GSR = "ENABLED";
    FD1P3AX array_255___i1834 (.D(array_0__7__N_2265[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[26] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1834.GSR = "ENABLED";
    FD1P3AX array_255___i1835 (.D(array_0__7__N_2265[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[26] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1835.GSR = "ENABLED";
    FD1P3AX array_255___i1836 (.D(array_0__7__N_2265[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[26] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1836.GSR = "ENABLED";
    FD1P3AX array_255___i1837 (.D(array_0__7__N_2265[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[26] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1837.GSR = "ENABLED";
    FD1P3AX array_255___i1838 (.D(array_0__7__N_2265[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[26] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1838.GSR = "ENABLED";
    FD1P3AX array_255___i1839 (.D(array_0__7__N_2265[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[26] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1839.GSR = "ENABLED";
    FD1P3AX array_255___i1840 (.D(array_0__7__N_2265[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[26] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1840.GSR = "ENABLED";
    FD1P3AX array_255___i1841 (.D(array_0__7__N_2257[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[25] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1841.GSR = "ENABLED";
    FD1P3AX array_255___i1842 (.D(array_0__7__N_2257[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[25] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1842.GSR = "ENABLED";
    FD1P3AX array_255___i1843 (.D(array_0__7__N_2257[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[25] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1843.GSR = "ENABLED";
    FD1P3AX array_255___i1844 (.D(array_0__7__N_2257[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[25] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1844.GSR = "ENABLED";
    FD1P3AX array_255___i1845 (.D(array_0__7__N_2257[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[25] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1845.GSR = "ENABLED";
    FD1P3AX array_255___i1846 (.D(array_0__7__N_2257[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[25] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1846.GSR = "ENABLED";
    FD1P3AX array_255___i1847 (.D(array_0__7__N_2257[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[25] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1847.GSR = "ENABLED";
    FD1P3AX array_255___i1848 (.D(array_0__7__N_2257[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[25] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1848.GSR = "ENABLED";
    FD1P3AX array_255___i1849 (.D(array_0__7__N_2249[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[24] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1849.GSR = "ENABLED";
    FD1P3AX array_255___i1850 (.D(array_0__7__N_2249[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[24] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1850.GSR = "ENABLED";
    FD1P3AX array_255___i1851 (.D(array_0__7__N_2249[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[24] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1851.GSR = "ENABLED";
    FD1P3AX array_255___i1852 (.D(array_0__7__N_2249[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[24] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1852.GSR = "ENABLED";
    FD1P3AX array_255___i1853 (.D(array_0__7__N_2249[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[24] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1853.GSR = "ENABLED";
    FD1P3AX array_255___i1854 (.D(array_0__7__N_2249[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[24] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1854.GSR = "ENABLED";
    FD1P3AX array_255___i1855 (.D(array_0__7__N_2249[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[24] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1855.GSR = "ENABLED";
    FD1P3AX array_255___i1856 (.D(array_0__7__N_2249[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[24] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1856.GSR = "ENABLED";
    FD1P3AX array_255___i1857 (.D(array_0__7__N_2241[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[23] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1857.GSR = "ENABLED";
    FD1P3AX array_255___i1858 (.D(array_0__7__N_2241[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[23] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1858.GSR = "ENABLED";
    FD1P3AX array_255___i1859 (.D(array_0__7__N_2241[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[23] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1859.GSR = "ENABLED";
    FD1P3AX array_255___i1860 (.D(array_0__7__N_2241[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[23] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1860.GSR = "ENABLED";
    FD1P3AX array_255___i1861 (.D(array_0__7__N_2241[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[23] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1861.GSR = "ENABLED";
    FD1P3AX array_255___i1862 (.D(array_0__7__N_2241[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[23] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1862.GSR = "ENABLED";
    FD1P3AX array_255___i1863 (.D(array_0__7__N_2241[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[23] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1863.GSR = "ENABLED";
    FD1P3AX array_255___i1864 (.D(array_0__7__N_2241[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[23] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1864.GSR = "ENABLED";
    FD1P3AX array_255___i1865 (.D(array_0__7__N_2233[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[22] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1865.GSR = "ENABLED";
    FD1P3AX array_255___i1866 (.D(array_0__7__N_2233[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[22] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1866.GSR = "ENABLED";
    FD1P3AX array_255___i1867 (.D(array_0__7__N_2233[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[22] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1867.GSR = "ENABLED";
    FD1P3AX array_255___i1868 (.D(array_0__7__N_2233[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[22] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1868.GSR = "ENABLED";
    FD1P3AX array_255___i1869 (.D(array_0__7__N_2233[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[22] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1869.GSR = "ENABLED";
    FD1P3AX array_255___i1870 (.D(array_0__7__N_2233[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[22] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1870.GSR = "ENABLED";
    FD1P3AX array_255___i1871 (.D(array_0__7__N_2233[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[22] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1871.GSR = "ENABLED";
    FD1P3AX array_255___i1872 (.D(array_0__7__N_2233[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[22] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1872.GSR = "ENABLED";
    FD1P3AX array_255___i1873 (.D(array_0__7__N_2225[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[21] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1873.GSR = "ENABLED";
    FD1P3AX array_255___i1874 (.D(array_0__7__N_2225[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[21] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1874.GSR = "ENABLED";
    FD1P3AX array_255___i1875 (.D(array_0__7__N_2225[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[21] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1875.GSR = "ENABLED";
    FD1P3AX array_255___i1876 (.D(array_0__7__N_2225[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[21] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1876.GSR = "ENABLED";
    FD1P3AX array_255___i1877 (.D(array_0__7__N_2225[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[21] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1877.GSR = "ENABLED";
    FD1P3AX array_255___i1878 (.D(array_0__7__N_2225[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[21] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1878.GSR = "ENABLED";
    FD1P3AX array_255___i1879 (.D(array_0__7__N_2225[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[21] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1879.GSR = "ENABLED";
    FD1P3AX array_255___i1880 (.D(array_0__7__N_2225[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[21] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1880.GSR = "ENABLED";
    FD1P3AX array_255___i1881 (.D(array_0__7__N_2217[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[20] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1881.GSR = "ENABLED";
    FD1P3AX array_255___i1882 (.D(array_0__7__N_2217[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[20] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1882.GSR = "ENABLED";
    FD1P3AX array_255___i1883 (.D(array_0__7__N_2217[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[20] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1883.GSR = "ENABLED";
    FD1P3AX array_255___i1884 (.D(array_0__7__N_2217[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[20] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1884.GSR = "ENABLED";
    FD1P3AX array_255___i1885 (.D(array_0__7__N_2217[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[20] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1885.GSR = "ENABLED";
    FD1P3AX array_255___i1886 (.D(array_0__7__N_2217[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[20] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1886.GSR = "ENABLED";
    FD1P3AX array_255___i1887 (.D(array_0__7__N_2217[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[20] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1887.GSR = "ENABLED";
    FD1P3AX array_255___i1888 (.D(array_0__7__N_2217[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[20] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1888.GSR = "ENABLED";
    FD1P3AX array_255___i1889 (.D(array_0__7__N_2209[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[19] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1889.GSR = "ENABLED";
    FD1P3AX array_255___i1890 (.D(array_0__7__N_2209[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[19] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1890.GSR = "ENABLED";
    FD1P3AX array_255___i1891 (.D(array_0__7__N_2209[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[19] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1891.GSR = "ENABLED";
    FD1P3AX array_255___i1892 (.D(array_0__7__N_2209[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[19] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1892.GSR = "ENABLED";
    FD1P3AX array_255___i1893 (.D(array_0__7__N_2209[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[19] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1893.GSR = "ENABLED";
    FD1P3AX array_255___i1894 (.D(array_0__7__N_2209[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[19] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1894.GSR = "ENABLED";
    FD1P3AX array_255___i1895 (.D(array_0__7__N_2209[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[19] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1895.GSR = "ENABLED";
    FD1P3AX array_255___i1896 (.D(array_0__7__N_2209[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[19] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1896.GSR = "ENABLED";
    FD1P3AX array_255___i1897 (.D(array_0__7__N_2201[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[18] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1897.GSR = "ENABLED";
    FD1P3AX array_255___i1898 (.D(array_0__7__N_2201[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[18] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1898.GSR = "ENABLED";
    FD1P3AX array_255___i1899 (.D(array_0__7__N_2201[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[18] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1899.GSR = "ENABLED";
    FD1P3AX array_255___i1900 (.D(array_0__7__N_2201[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[18] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1900.GSR = "ENABLED";
    FD1P3AX array_255___i1901 (.D(array_0__7__N_2201[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[18] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1901.GSR = "ENABLED";
    FD1P3AX array_255___i1902 (.D(array_0__7__N_2201[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[18] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1902.GSR = "ENABLED";
    FD1P3AX array_255___i1903 (.D(array_0__7__N_2201[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[18] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1903.GSR = "ENABLED";
    FD1P3AX array_255___i1904 (.D(array_0__7__N_2201[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[18] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1904.GSR = "ENABLED";
    FD1P3AX array_255___i1905 (.D(array_0__7__N_2193[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[17] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1905.GSR = "ENABLED";
    FD1P3AX array_255___i1906 (.D(array_0__7__N_2193[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[17] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1906.GSR = "ENABLED";
    FD1P3AX array_255___i1907 (.D(array_0__7__N_2193[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[17] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1907.GSR = "ENABLED";
    FD1P3AX array_255___i1908 (.D(array_0__7__N_2193[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[17] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1908.GSR = "ENABLED";
    FD1P3AX array_255___i1909 (.D(array_0__7__N_2193[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[17] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1909.GSR = "ENABLED";
    FD1P3AX array_255___i1910 (.D(array_0__7__N_2193[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[17] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1910.GSR = "ENABLED";
    FD1P3AX array_255___i1911 (.D(array_0__7__N_2193[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[17] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1911.GSR = "ENABLED";
    FD1P3AX array_255___i1912 (.D(array_0__7__N_2193[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[17] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1912.GSR = "ENABLED";
    FD1P3AX array_255___i1913 (.D(array_0__7__N_2185[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[16] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1913.GSR = "ENABLED";
    FD1P3AX array_255___i1914 (.D(array_0__7__N_2185[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[16] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1914.GSR = "ENABLED";
    FD1P3AX array_255___i1915 (.D(array_0__7__N_2185[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[16] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1915.GSR = "ENABLED";
    FD1P3AX array_255___i1916 (.D(array_0__7__N_2185[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[16] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1916.GSR = "ENABLED";
    FD1P3AX array_255___i1917 (.D(array_0__7__N_2185[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[16] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1917.GSR = "ENABLED";
    FD1P3AX array_255___i1918 (.D(array_0__7__N_2185[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[16] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1918.GSR = "ENABLED";
    FD1P3AX array_255___i1919 (.D(array_0__7__N_2185[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[16] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1919.GSR = "ENABLED";
    FD1P3AX array_255___i1920 (.D(array_0__7__N_2185[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[16] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1920.GSR = "ENABLED";
    FD1P3AX array_255___i1921 (.D(array_0__7__N_2177[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[15] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1921.GSR = "ENABLED";
    FD1P3AX array_255___i1922 (.D(array_0__7__N_2177[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[15] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1922.GSR = "ENABLED";
    FD1P3AX array_255___i1923 (.D(array_0__7__N_2177[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[15] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1923.GSR = "ENABLED";
    FD1P3AX array_255___i1924 (.D(array_0__7__N_2177[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[15] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1924.GSR = "ENABLED";
    FD1P3AX array_255___i1925 (.D(array_0__7__N_2177[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[15] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1925.GSR = "ENABLED";
    FD1P3AX array_255___i1926 (.D(array_0__7__N_2177[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[15] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1926.GSR = "ENABLED";
    FD1P3AX array_255___i1927 (.D(array_0__7__N_2177[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[15] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1927.GSR = "ENABLED";
    FD1P3AX array_255___i1928 (.D(array_0__7__N_2177[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[15] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1928.GSR = "ENABLED";
    FD1P3AX array_255___i1929 (.D(array_0__7__N_2169[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[14] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1929.GSR = "ENABLED";
    FD1P3AX array_255___i1930 (.D(array_0__7__N_2169[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[14] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1930.GSR = "ENABLED";
    FD1P3AX array_255___i1931 (.D(array_0__7__N_2169[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[14] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1931.GSR = "ENABLED";
    FD1P3AX array_255___i1932 (.D(array_0__7__N_2169[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[14] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1932.GSR = "ENABLED";
    FD1P3AX array_255___i1933 (.D(array_0__7__N_2169[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[14] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1933.GSR = "ENABLED";
    FD1P3AX array_255___i1934 (.D(array_0__7__N_2169[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[14] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1934.GSR = "ENABLED";
    FD1P3AX array_255___i1935 (.D(array_0__7__N_2169[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[14] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1935.GSR = "ENABLED";
    FD1P3AX array_255___i1936 (.D(array_0__7__N_2169[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[14] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1936.GSR = "ENABLED";
    FD1P3AX array_255___i1937 (.D(array_0__7__N_2161[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[13] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1937.GSR = "ENABLED";
    FD1P3AX array_255___i1938 (.D(array_0__7__N_2161[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[13] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1938.GSR = "ENABLED";
    FD1P3AX array_255___i1939 (.D(array_0__7__N_2161[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[13] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1939.GSR = "ENABLED";
    FD1P3AX array_255___i1940 (.D(array_0__7__N_2161[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[13] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1940.GSR = "ENABLED";
    FD1P3AX array_255___i1941 (.D(array_0__7__N_2161[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[13] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1941.GSR = "ENABLED";
    FD1P3AX array_255___i1942 (.D(array_0__7__N_2161[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[13] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1942.GSR = "ENABLED";
    FD1P3AX array_255___i1943 (.D(array_0__7__N_2161[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[13] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1943.GSR = "ENABLED";
    FD1P3AX array_255___i1944 (.D(array_0__7__N_2161[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[13] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1944.GSR = "ENABLED";
    FD1P3AX array_255___i1945 (.D(array_0__7__N_2153[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[12] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1945.GSR = "ENABLED";
    FD1P3AX array_255___i1946 (.D(array_0__7__N_2153[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[12] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1946.GSR = "ENABLED";
    FD1P3AX array_255___i1947 (.D(array_0__7__N_2153[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[12] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1947.GSR = "ENABLED";
    FD1P3AX array_255___i1948 (.D(array_0__7__N_2153[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[12] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1948.GSR = "ENABLED";
    FD1P3AX array_255___i1949 (.D(array_0__7__N_2153[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[12] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1949.GSR = "ENABLED";
    FD1P3AX array_255___i1950 (.D(array_0__7__N_2153[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[12] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1950.GSR = "ENABLED";
    FD1P3AX array_255___i1951 (.D(array_0__7__N_2153[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[12] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1951.GSR = "ENABLED";
    FD1P3AX array_255___i1952 (.D(array_0__7__N_2153[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[12] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1952.GSR = "ENABLED";
    FD1P3AX array_255___i1953 (.D(array_0__7__N_2145[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[11] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1953.GSR = "ENABLED";
    FD1P3AX array_255___i1954 (.D(array_0__7__N_2145[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[11] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1954.GSR = "ENABLED";
    FD1P3AX array_255___i1955 (.D(array_0__7__N_2145[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[11] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1955.GSR = "ENABLED";
    FD1P3AX array_255___i1956 (.D(array_0__7__N_2145[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[11] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1956.GSR = "ENABLED";
    FD1P3AX array_255___i1957 (.D(array_0__7__N_2145[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[11] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1957.GSR = "ENABLED";
    FD1P3AX array_255___i1958 (.D(array_0__7__N_2145[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[11] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1958.GSR = "ENABLED";
    FD1P3AX array_255___i1959 (.D(array_0__7__N_2145[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[11] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1959.GSR = "ENABLED";
    FD1P3AX array_255___i1960 (.D(array_0__7__N_2145[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[11] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1960.GSR = "ENABLED";
    FD1P3AX array_255___i1961 (.D(array_0__7__N_2137[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[10] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1961.GSR = "ENABLED";
    FD1P3AX array_255___i1962 (.D(array_0__7__N_2137[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[10] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1962.GSR = "ENABLED";
    FD1P3AX array_255___i1963 (.D(array_0__7__N_2137[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[10] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1963.GSR = "ENABLED";
    FD1P3AX array_255___i1964 (.D(array_0__7__N_2137[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[10] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1964.GSR = "ENABLED";
    FD1P3AX array_255___i1965 (.D(array_0__7__N_2137[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[10] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1965.GSR = "ENABLED";
    FD1P3AX array_255___i1966 (.D(array_0__7__N_2137[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[10] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1966.GSR = "ENABLED";
    FD1P3AX array_255___i1967 (.D(array_0__7__N_2137[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[10] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1967.GSR = "ENABLED";
    FD1P3AX array_255___i1968 (.D(array_0__7__N_2137[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[10] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1968.GSR = "ENABLED";
    FD1P3AX array_255___i1969 (.D(array_0__7__N_2129[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[9] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1969.GSR = "ENABLED";
    FD1P3AX array_255___i1970 (.D(array_0__7__N_2129[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[9] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1970.GSR = "ENABLED";
    FD1P3AX array_255___i1971 (.D(array_0__7__N_2129[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[9] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1971.GSR = "ENABLED";
    FD1P3AX array_255___i1972 (.D(array_0__7__N_2129[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[9] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1972.GSR = "ENABLED";
    FD1P3AX array_255___i1973 (.D(array_0__7__N_2129[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[9] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1973.GSR = "ENABLED";
    FD1P3AX array_255___i1974 (.D(array_0__7__N_2129[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[9] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1974.GSR = "ENABLED";
    FD1P3AX array_255___i1975 (.D(array_0__7__N_2129[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[9] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1975.GSR = "ENABLED";
    FD1P3AX array_255___i1976 (.D(array_0__7__N_2129[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[9] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1976.GSR = "ENABLED";
    FD1P3AX array_255___i1977 (.D(array_0__7__N_2121[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[8] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1977.GSR = "ENABLED";
    FD1P3AX array_255___i1978 (.D(array_0__7__N_2121[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[8] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1978.GSR = "ENABLED";
    FD1P3AX array_255___i1979 (.D(array_0__7__N_2121[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[8] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1979.GSR = "ENABLED";
    FD1P3AX array_255___i1980 (.D(array_0__7__N_2121[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[8] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1980.GSR = "ENABLED";
    FD1P3AX array_255___i1981 (.D(array_0__7__N_2121[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[8] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1981.GSR = "ENABLED";
    FD1P3AX array_255___i1982 (.D(array_0__7__N_2121[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[8] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1982.GSR = "ENABLED";
    FD1P3AX array_255___i1983 (.D(array_0__7__N_2121[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[8] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1983.GSR = "ENABLED";
    FD1P3AX array_255___i1984 (.D(array_0__7__N_2121[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[8] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1984.GSR = "ENABLED";
    FD1P3AX array_255___i1985 (.D(array_0__7__N_2113[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[7] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1985.GSR = "ENABLED";
    FD1P3AX array_255___i1986 (.D(array_0__7__N_2113[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[7] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1986.GSR = "ENABLED";
    FD1P3AX array_255___i1987 (.D(array_0__7__N_2113[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[7] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1987.GSR = "ENABLED";
    FD1P3AX array_255___i1988 (.D(array_0__7__N_2113[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[7] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1988.GSR = "ENABLED";
    FD1P3AX array_255___i1989 (.D(array_0__7__N_2113[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[7] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1989.GSR = "ENABLED";
    FD1P3AX array_255___i1990 (.D(array_0__7__N_2113[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[7] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1990.GSR = "ENABLED";
    FD1P3AX array_255___i1991 (.D(array_0__7__N_2113[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[7] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1991.GSR = "ENABLED";
    FD1P3AX array_255___i1992 (.D(array_0__7__N_2113[7]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[7] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1992.GSR = "ENABLED";
    FD1P3AX array_255___i1993 (.D(array_0__7__N_2105[0]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[6] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1993.GSR = "ENABLED";
    FD1P3AX array_255___i1994 (.D(array_0__7__N_2105[1]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[6] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1994.GSR = "ENABLED";
    FD1P3AX array_255___i1995 (.D(array_0__7__N_2105[2]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[6] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1995.GSR = "ENABLED";
    FD1P3AX array_255___i1996 (.D(array_0__7__N_2105[3]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[6] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1996.GSR = "ENABLED";
    FD1P3AX array_255___i1997 (.D(array_0__7__N_2105[4]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[6] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1997.GSR = "ENABLED";
    FD1P3AX array_255___i1998 (.D(array_0__7__N_2105[5]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[6] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1998.GSR = "ENABLED";
    FD1P3AX array_255___i1999 (.D(array_0__7__N_2105[6]), .SP(clk_c_enable_2007), 
            .CK(clk_c), .Q(\array[6] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i1999.GSR = "ENABLED";
    FD1P3AX array_255___i2000 (.D(array_0__7__N_2105[7]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[6] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2000.GSR = "ENABLED";
    FD1P3AX array_255___i2001 (.D(array_0__7__N_2097[0]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[5] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2001.GSR = "ENABLED";
    FD1P3AX array_255___i2002 (.D(array_0__7__N_2097[1]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[5] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2002.GSR = "ENABLED";
    FD1P3AX array_255___i2003 (.D(array_0__7__N_2097[2]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[5] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2003.GSR = "ENABLED";
    FD1P3AX array_255___i2004 (.D(array_0__7__N_2097[3]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[5] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2004.GSR = "ENABLED";
    FD1P3AX array_255___i2005 (.D(array_0__7__N_2097[4]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[5] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2005.GSR = "ENABLED";
    FD1P3AX array_255___i2006 (.D(array_0__7__N_2097[5]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[5] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2006.GSR = "ENABLED";
    FD1P3AX array_255___i2007 (.D(array_0__7__N_2097[6]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[5] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2007.GSR = "ENABLED";
    FD1P3AX array_255___i2008 (.D(array_0__7__N_2097[7]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[5] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2008.GSR = "ENABLED";
    FD1P3AX array_255___i2009 (.D(array_0__7__N_2089[0]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[4] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2009.GSR = "ENABLED";
    FD1P3AX array_255___i2010 (.D(array_0__7__N_2089[1]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[4] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2010.GSR = "ENABLED";
    FD1P3AX array_255___i2011 (.D(array_0__7__N_2089[2]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[4] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2011.GSR = "ENABLED";
    FD1P3AX array_255___i2012 (.D(array_0__7__N_2089[3]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[4] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2012.GSR = "ENABLED";
    FD1P3AX array_255___i2013 (.D(array_0__7__N_2089[4]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[4] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2013.GSR = "ENABLED";
    FD1P3AX array_255___i2014 (.D(array_0__7__N_2089[5]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[4] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2014.GSR = "ENABLED";
    FD1P3AX array_255___i2015 (.D(array_0__7__N_2089[6]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[4] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2015.GSR = "ENABLED";
    FD1P3AX array_255___i2016 (.D(array_0__7__N_2089[7]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[4] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2016.GSR = "ENABLED";
    FD1P3AX array_255___i2017 (.D(array_0__7__N_2081[0]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[3] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2017.GSR = "ENABLED";
    FD1P3AX array_255___i2018 (.D(array_0__7__N_2081[1]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[3] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2018.GSR = "ENABLED";
    FD1P3AX array_255___i2019 (.D(array_0__7__N_2081[2]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[3] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2019.GSR = "ENABLED";
    FD1P3AX array_255___i2020 (.D(array_0__7__N_2081[3]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[3] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2020.GSR = "ENABLED";
    FD1P3AX array_255___i2021 (.D(array_0__7__N_2081[4]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[3] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2021.GSR = "ENABLED";
    FD1P3AX array_255___i2022 (.D(array_0__7__N_2081[5]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[3] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2022.GSR = "ENABLED";
    FD1P3AX array_255___i2023 (.D(array_0__7__N_2081[6]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[3] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2023.GSR = "ENABLED";
    FD1P3AX array_255___i2024 (.D(array_0__7__N_2081[7]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[3] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2024.GSR = "ENABLED";
    FD1P3AX array_255___i2025 (.D(array_0__7__N_2073[0]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[2] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2025.GSR = "ENABLED";
    FD1P3AX array_255___i2026 (.D(array_0__7__N_2073[1]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[2] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2026.GSR = "ENABLED";
    FD1P3AX array_255___i2027 (.D(array_0__7__N_2073[2]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[2] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2027.GSR = "ENABLED";
    FD1P3AX array_255___i2028 (.D(array_0__7__N_2073[3]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[2] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2028.GSR = "ENABLED";
    FD1P3AX array_255___i2029 (.D(array_0__7__N_2073[4]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[2] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2029.GSR = "ENABLED";
    FD1P3AX array_255___i2030 (.D(array_0__7__N_2073[5]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[2] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2030.GSR = "ENABLED";
    FD1P3AX array_255___i2031 (.D(array_0__7__N_2073[6]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[2] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2031.GSR = "ENABLED";
    FD1P3AX array_255___i2032 (.D(array_0__7__N_2073[7]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[2] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2032.GSR = "ENABLED";
    FD1P3AX array_255___i2033 (.D(array_0__7__N_2065[0]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[1] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2033.GSR = "ENABLED";
    FD1P3AX array_255___i2034 (.D(array_0__7__N_2065[1]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[1] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2034.GSR = "ENABLED";
    FD1P3AX array_255___i2035 (.D(array_0__7__N_2065[2]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[1] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2035.GSR = "ENABLED";
    FD1P3AX array_255___i2036 (.D(array_0__7__N_2065[3]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[1] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2036.GSR = "ENABLED";
    FD1P3AX array_255___i2037 (.D(array_0__7__N_2065[4]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[1] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2037.GSR = "ENABLED";
    FD1P3AX array_255___i2038 (.D(array_0__7__N_2065[5]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[1] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2038.GSR = "ENABLED";
    FD1P3AX array_255___i2039 (.D(array_0__7__N_2065[6]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[1] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2039.GSR = "ENABLED";
    FD1P3AX array_255___i2040 (.D(array_0__7__N_2065[7]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[1] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2040.GSR = "ENABLED";
    FD1P3AX array_255___i2041 (.D(array_0__7__N_2057[0]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[0] [0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2041.GSR = "ENABLED";
    FD1P3AX array_255___i2042 (.D(array_0__7__N_2057[1]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[0] [1]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2042.GSR = "ENABLED";
    FD1P3AX array_255___i2043 (.D(array_0__7__N_2057[2]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[0] [2]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2043.GSR = "ENABLED";
    FD1P3AX array_255___i2044 (.D(array_0__7__N_2057[3]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[0] [3]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2044.GSR = "ENABLED";
    FD1P3AX array_255___i2045 (.D(array_0__7__N_2057[4]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[0] [4]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2045.GSR = "ENABLED";
    FD1P3AX array_255___i2046 (.D(array_0__7__N_2057[5]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[0] [5]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2046.GSR = "ENABLED";
    FD1P3AX array_255___i2047 (.D(array_0__7__N_2057[6]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[0] [6]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2047.GSR = "ENABLED";
    FD1P3AX array_255___i2048 (.D(array_0__7__N_2057[7]), .SP(clk_c_enable_2056), 
            .CK(clk_c), .Q(\array[0] [7]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam array_255___i2048.GSR = "ENABLED";
    FD1P3AX r_addr_i0_i0 (.D(addr_c_0), .SP(clk_c_enable_2057), .CK(clk_c), 
            .Q(r_addr[0]));   // c:/users/user/documents/fpga/srdydrdy_lib/trunk/rtl/verilog/memory/behave1p_mem.v(27[10] 37[8])
    defparam r_addr_i0_i0.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

